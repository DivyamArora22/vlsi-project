VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LAYER contactResistance REAL ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MANUFACTURINGGRID 0.0025 ;
LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER poly
  TYPE MASTERSLICE ;
END poly

LAYER contact
  TYPE CUT ;
  SPACING 0.075 ;
  PROPERTY contactResistance 10.5 ;
END contact

LAYER metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 0.19 ;
  WIDTH 0.065 ;
  SPACING 0.065 ;
  SPACING 0.065 SAMENET ;
  RESISTANCE RPERSQ 0.38 ;
END metal1

LAYER via1
  TYPE CUT ;
  SPACING 0.075 ;
  WIDTH 0.065 ;
  PROPERTY contactResistance 5.69 ;
END via1

LAYER metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.19 0.19 ;
  WIDTH 0.07 ;
  SPACING 0.075 ;
  SPACING 0.07 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal2

LAYER via2
  TYPE CUT ;
  SPACING 0.085 ;
  WIDTH 0.07 ;
  PROPERTY contactResistance 11.39 ;
END via2

LAYER metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.19 0.19 ;
  WIDTH 0.07 ;
  SPACING 0.07 ;
  SPACING 0.07 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal3

LAYER via3
  TYPE CUT ;
  SPACING 0.085 ;
  WIDTH 0.07 ;
  PROPERTY contactResistance 16.73 ;
END via3

LAYER metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.285 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  SPACING 0.14 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal4

LAYER via4
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  PROPERTY contactResistance 21.44 ;
END via4

LAYER metal5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.285 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  SPACING 0.14 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal5

LAYER via5
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  PROPERTY contactResistance 24.08 ;
END via5

LAYER metal6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.285 0.285 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  SPACING 0.14 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal6

LAYER via6
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  PROPERTY contactResistance 11.39 ;
END via6

LAYER metal7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.855 0.855 ;
  WIDTH 0.4 ;
  SPACING 0.44 ;
  SPACING 0.44 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal7

LAYER via7
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  PROPERTY contactResistance 5.69 ;
END via7

LAYER metal8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.855 0.855 ;
  WIDTH 0.4 ;
  SPACING 0.44 ;
  SPACING 0.44 SAMENET ;
  RESISTANCE RPERSQ 0.25 ;
END metal8

LAYER via8
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  PROPERTY contactResistance 16.73 ;
END via8

LAYER metal9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.71 1.71 ;
  WIDTH 0.8 ;
  SPACING 0.8 ;
  SPACING 0.8 SAMENET ;
  RESISTANCE RPERSQ 0.21 ;
END metal9

LAYER via9
  TYPE CUT ;
  SPACING 0.88 ;
  WIDTH 0.8 ;
  PROPERTY contactResistance 21.44 ;
END via9

LAYER metal10
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.71 1.71 ;
  WIDTH 0.4 ;
  SPACING 0.8 ;
  SPACING 0.8 SAMENET ;
  RESISTANCE RPERSQ 0.21 ;
END metal10

VIARULE M2_M1 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
    SPACING 0.14 BY 0.14 ;
END M2_M1

VIARULE M3_M2 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END M3_M2

VIARULE M4_M3 GENERATE
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.155 BY 0.155 ;
END M4_M3

VIARULE M5_M4 GENERATE
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M5_M4

VIARULE M6_M5 GENERATE
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M6_M5

VIARULE M7_M6 GENERATE
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER metal7 ;
    ENCLOSURE 0.13 0.13 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END M7_M6

VIARULE M8_M7 GENERATE
  LAYER metal7 ;
    ENCLOSURE 0 0 ;
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.8 BY 0.8 ;
END M8_M7

VIARULE M9_M8 GENERATE
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER metal9 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.8 BY 0.8 ;
END M9_M8

VIARULE M10_M9 GENERATE
  LAYER metal9 ;
    ENCLOSURE 0 0 ;
  LAYER metal10 ;
    ENCLOSURE 0 0 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 1.6 BY 1.6 ;
END M10_M9

VIARULE M1_POLY GENERATE
  LAYER poly ;
    ENCLOSURE 0 0 ;
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
  LAYER contact ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
    SPACING 0.14 BY 0.14 ;
END M1_POLY

VIA M2_M1_via DEFAULT
  LAYER metal1 ;
    RECT -0.0675 -0.0325 0.0675 0.0325 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.035 -0.0675 0.035 0.0675 ;
END M2_M1_via

VIA M3_M2_via DEFAULT
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END M3_M2_via

VIA M4_M3_via DEFAULT
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M4_M3_via

VIA M5_M4_via DEFAULT
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M5_M4_via

VIA M6_M5_via DEFAULT
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M6_M5_via

VIA M7_M6_via DEFAULT
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END M7_M6_via

VIA M8_M7_via DEFAULT
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END M8_M7_via

VIA M9_M8_via DEFAULT
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END M9_M8_via

VIA M10_M9_via DEFAULT
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER metal10 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END M10_M9_via

VIA M2_M1_viaB DEFAULT
  LAYER metal1 ;
    RECT -0.0675 -0.0325 0.0675 0.0325 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.0675 -0.035 0.0675 0.035 ;
END M2_M1_viaB

VIA M2_M1_viaC DEFAULT
  LAYER metal1 ;
    RECT -0.0325 -0.0675 0.0325 0.0675 ;
  LAYER via1 ;
    RECT -0.0325 -0.0325 0.0325 0.0325 ;
  LAYER metal2 ;
    RECT -0.035 -0.0675 0.035 0.0675 ;
END M2_M1_viaC

VIA M3_M2_viaB DEFAULT
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END M3_M2_viaB

VIA M3_M2_viaC DEFAULT
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END M3_M2_viaC

VIA M4_M3_viaB DEFAULT
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END M4_M3_viaB

SITE CoreSite
  CLASS CORE ;
  SIZE 0.005 BY 1.45 ;
END CoreSite

MACRO and2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN and2 0 0.1 ;
  SIZE 0.8025 BY 1.45 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.45 0.8025 1.65 ;
        RECT 0.6775 1.2375 0.7425 1.65 ;
        RECT 0.3025 1.26 0.3675 1.65 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.8025 0.2 ;
        RECT 0.3025 0 0.3675 0.4225 ;
    END
  END vss!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.335 0.6025 0.4 0.7375 ;
      LAYER metal2 ;
        RECT 0.3325 0.6025 0.4025 0.7375 ;
      LAYER via1 ;
        RECT 0.335 0.6375 0.4 0.7025 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.545 0.8925 0.61 1.0275 ;
      LAYER metal2 ;
        RECT 0.5425 0.8925 0.6125 1.0275 ;
      LAYER via1 ;
        RECT 0.545 0.9275 0.61 0.9925 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.275 0.125 1.3725 ;
        RECT 0.0575 0.79 0.125 0.925 ;
      LAYER metal2 ;
        RECT 0.055 0.79 0.125 0.925 ;
      LAYER via1 ;
        RECT 0.0575 0.825 0.1225 0.89 ;
    END
  END Y
  OBS
    LAYER metal1 ;
      RECT 0.49 1.0925 0.555 1.36 ;
      RECT 0.2125 1.095 0.555 1.16 ;
      RECT 0.685 0.3475 0.75 1.1575 ;
      RECT 0.49 1.0925 0.75 1.1575 ;
      RECT 0.19 1.0225 0.255 1.1575 ;
      RECT 0.6775 0.315 0.7425 0.45 ;
  END
END and2

MACRO aoi21
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN aoi21 0 0.1 ;
  SIZE 0.75 BY 1.45 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.45 0.75 1.65 ;
        RECT 0.06 1.0375 0.125 1.65 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.75 0.2 ;
        RECT 0.625 0 0.69 0.36 ;
        RECT 0.06 0 0.125 0.4125 ;
    END
  END vss!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.255 0.86 0.39 0.925 ;
      LAYER metal2 ;
        RECT 0.255 0.8575 0.39 0.9275 ;
      LAYER via1 ;
        RECT 0.29 0.86 0.355 0.925 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.48 0.7825 0.545 0.9175 ;
      LAYER metal2 ;
        RECT 0.4775 0.7825 0.5475 0.9175 ;
      LAYER via1 ;
        RECT 0.48 0.8175 0.545 0.8825 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.08 0.825 0.145 0.96 ;
      LAYER metal2 ;
        RECT 0.0775 0.825 0.1475 0.96 ;
      LAYER via1 ;
        RECT 0.08 0.86 0.145 0.925 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6375 0.79 0.7125 0.925 ;
        RECT 0.4375 1.0025 0.7025 1.0675 ;
        RECT 0.6375 0.575 0.7025 1.0675 ;
        RECT 0.2475 0.575 0.7025 0.64 ;
        RECT 0.4375 1.0025 0.5025 1.2175 ;
        RECT 0.2475 0.265 0.3125 0.64 ;
      LAYER metal2 ;
        RECT 0.645 0.79 0.715 0.925 ;
      LAYER via1 ;
        RECT 0.6475 0.825 0.7125 0.89 ;
    END
  END Y
  OBS
    LAYER metal1 ;
      RECT 0.625 1.1325 0.69 1.2725 ;
      RECT 0.2475 1.135 0.3125 1.275 ;
    LAYER metal2 ;
      RECT 0.245 1 0.315 1.275 ;
      RECT 0.6225 1 0.6925 1.2725 ;
      RECT 0.245 1 0.6925 1.07 ;
    LAYER via1 ;
      RECT 0.625 1.1725 0.69 1.2375 ;
      RECT 0.2475 1.175 0.3125 1.24 ;
  END
END aoi21

MACRO buf
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN buf 0 0.1 ;
  SIZE 0.605 BY 1.45 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.45 0.605 1.65 ;
        RECT 0.27 1.23 0.335 1.65 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.605 0.2 ;
        RECT 0.27 0 0.335 0.44 ;
    END
  END vss!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3225 0.7 0.3875 0.835 ;
      LAYER metal2 ;
        RECT 0.32 0.7 0.39 0.835 ;
      LAYER via1 ;
        RECT 0.3225 0.735 0.3875 0.8 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.08 0.27 0.145 1.3725 ;
        RECT 0.0375 0.535 0.145 0.67 ;
      LAYER metal2 ;
        RECT 0.035 0.535 0.105 0.67 ;
      LAYER via1 ;
        RECT 0.0375 0.57 0.1025 0.635 ;
    END
  END Y
  OBS
    LAYER metal1 ;
      RECT 0.4575 0.265 0.5225 1.3725 ;
      RECT 0.4575 0.9725 0.5675 1.1075 ;
      RECT 0.21 0.9725 0.275 1.1075 ;
    LAYER metal2 ;
      RECT 0.5 0.9725 0.57 1.1075 ;
      RECT 0.2075 0.9725 0.2775 1.1075 ;
      RECT 0.2075 1.005 0.57 1.075 ;
    LAYER via1 ;
      RECT 0.5025 1.0075 0.5675 1.0725 ;
      RECT 0.21 1.0075 0.275 1.0725 ;
  END
END buf

MACRO dff
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN dff 0 0.1 ;
  SIZE 3.7025 BY 1.45 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.45 3.7 1.65 ;
        RECT 3.305 1.2475 3.37 1.65 ;
        RECT 1.9375 1.2475 2.0025 1.65 ;
        RECT 1.0025 1.22 1.0675 1.65 ;
        RECT 0.25 1.2 0.315 1.65 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 3.7025 0.2 ;
        RECT 3.305 0 3.37 0.385 ;
        RECT 1.9375 0 2.0025 0.385 ;
        RECT 1.0025 0 1.0675 0.385 ;
        RECT 0.25 0 0.315 0.385 ;
    END
  END vss!
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.295 0.6825 0.36 0.8175 ;
      LAYER metal2 ;
        RECT 0.2925 0.6825 0.3625 0.8175 ;
      LAYER via1 ;
        RECT 0.295 0.7175 0.36 0.7825 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.035 0.4525 1.1 0.5875 ;
      LAYER metal2 ;
        RECT 1.0325 0.4525 1.1025 0.5875 ;
      LAYER via1 ;
        RECT 1.035 0.4875 1.1 0.5525 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.655 0.265 0.72 1.3575 ;
      LAYER metal2 ;
        RECT 0.6525 1.0825 0.7225 1.2175 ;
      LAYER via1 ;
        RECT 0.655 1.1175 0.72 1.1825 ;
    END
  END Q
  OBS
    LAYER metal1 ;
      RECT 2.1775 0.265 2.2425 1.355 ;
      RECT 1.8425 0.99 1.9075 1.125 ;
      RECT 1.845 0.83 1.91 1.065 ;
      RECT 1.845 0.83 2.2425 0.895 ;
      RECT 1.4525 0.265 1.5175 1.3125 ;
      RECT 1.4525 1.1275 1.5475 1.2625 ;
      RECT 1.19 1.22 1.255 1.355 ;
      RECT 1.1875 0.265 1.2525 1.3525 ;
      RECT 1.1875 0.265 1.255 0.4 ;
      RECT 0.4375 0.265 0.5025 1.3475 ;
      RECT 0.4375 0.69 0.5625 0.825 ;
      RECT 0.0625 0.265 0.1275 1.345 ;
      RECT 0.06 1.2075 0.1275 1.3425 ;
      RECT 0.0625 0.8725 0.13 1.0075 ;
      RECT 0.06 0.265 0.1275 0.4 ;
      RECT 3.545 0.265 3.61 1.2925 ;
      RECT 3.405 1.03 3.47 1.165 ;
      RECT 3.21 1.03 3.275 1.165 ;
      RECT 2.9975 0.265 3.0625 1.3725 ;
      RECT 2.8575 0.405 2.9225 0.54 ;
      RECT 2.835 1.0225 2.9 1.1575 ;
      RECT 2.6425 0.265 2.7075 1.2925 ;
      RECT 2.3525 1.015 2.4175 1.15 ;
      RECT 2.3125 0.565 2.3775 0.7 ;
      RECT 2.0375 1.025 2.1025 1.16 ;
      RECT 1.7125 0.265 1.7775 1.3825 ;
      RECT 1.5825 0.565 1.6475 0.7 ;
      RECT 1.5825 0.9225 1.6475 1.0575 ;
      RECT 1.3225 0.405 1.3875 0.54 ;
      RECT 1.3225 1 1.3875 1.135 ;
      RECT 0.88 0.455 0.945 0.59 ;
      RECT 0.195 0.4525 0.26 0.5875 ;
    LAYER metal2 ;
      RECT 3.5425 0.265 3.6125 0.905 ;
      RECT 0.8775 0.455 0.9475 0.59 ;
      RECT 0.875 0.265 0.945 0.49 ;
      RECT 0.875 0.265 3.6125 0.335 ;
      RECT 3.2075 1.365 3.6125 1.435 ;
      RECT 3.5425 1.1575 3.6125 1.435 ;
      RECT 3.2075 1.03 3.2775 1.435 ;
      RECT 2.64 0.85 2.71 1.2925 ;
      RECT 3.4025 0.85 3.4725 1.165 ;
      RECT 2.64 0.85 3.4725 0.92 ;
      RECT 2.345 0.7825 2.415 1.155 ;
      RECT 2.345 1.015 2.42 1.15 ;
      RECT 1.58 0.7825 1.65 1.0575 ;
      RECT 1.58 0.7825 2.5225 0.8525 ;
      RECT 2.4525 0.425 2.5225 0.8525 ;
      RECT 0.495 0.67 0.565 0.825 ;
      RECT 0.4875 0.67 1.2425 0.74 ;
      RECT 1.1725 0.425 1.2425 0.74 ;
      RECT 2.855 0.405 2.925 0.54 ;
      RECT 1.32 0.405 1.39 0.54 ;
      RECT 1.1725 0.425 2.925 0.495 ;
      RECT 1.32 1.365 2.905 1.435 ;
      RECT 2.835 1.035 2.905 1.435 ;
      RECT 1.32 0.9 1.39 1.435 ;
      RECT 2.8325 1.0225 2.9025 1.1575 ;
      RECT 1.32 0.9 1.3975 1.135 ;
      RECT 1.3175 0.61 1.3875 1.1225 ;
      RECT 0.0625 0.8725 0.1325 1.0075 ;
      RECT 0.0625 0.9 1.3975 0.97 ;
      RECT 2.31 0.565 2.38 0.7 ;
      RECT 1.58 0.565 1.65 0.7 ;
      RECT 1.3175 0.61 2.38 0.68 ;
      RECT 1.48 1.1275 1.55 1.2625 ;
      RECT 1.48 1.1275 2.1025 1.1975 ;
      RECT 2.035 1.025 2.105 1.16 ;
      RECT 2.0325 1.0575 2.105 1.16 ;
      RECT 0.435 0.455 0.505 0.59 ;
      RECT 0.1925 0.4525 0.2625 0.5875 ;
      RECT 0.1875 0.4825 0.5075 0.5525 ;
    LAYER via1 ;
      RECT 3.545 0.805 3.61 0.87 ;
      RECT 3.545 1.1925 3.61 1.2575 ;
      RECT 3.405 1.065 3.47 1.13 ;
      RECT 3.21 1.065 3.275 1.13 ;
      RECT 2.8575 0.44 2.9225 0.505 ;
      RECT 2.835 1.0575 2.9 1.1225 ;
      RECT 2.6425 1.1925 2.7075 1.2575 ;
      RECT 2.3525 1.05 2.4175 1.115 ;
      RECT 2.3125 0.6 2.3775 0.665 ;
      RECT 2.0375 1.06 2.1025 1.125 ;
      RECT 1.5825 0.6 1.6475 0.665 ;
      RECT 1.5825 0.9575 1.6475 1.0225 ;
      RECT 1.4825 1.1625 1.5475 1.2275 ;
      RECT 1.3225 0.44 1.3875 0.505 ;
      RECT 1.3225 1.035 1.3875 1.1 ;
      RECT 0.88 0.49 0.945 0.555 ;
      RECT 0.4975 0.725 0.5625 0.79 ;
      RECT 0.4375 0.49 0.5025 0.555 ;
      RECT 0.195 0.4875 0.26 0.5525 ;
      RECT 0.065 0.9075 0.13 0.9725 ;
  END
END dff

MACRO inv
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN inv 0 0.1 ;
  SIZE 0.385 BY 1.45 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.45 0.385 1.65 ;
        RECT 0.06 1.23 0.125 1.65 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.385 0.2 ;
        RECT 0.06 0 0.125 0.415 ;
    END
  END vss!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.0925 0.825 0.1575 0.96 ;
      LAYER metal2 ;
        RECT 0.09 0.825 0.16 0.96 ;
      LAYER via1 ;
        RECT 0.0925 0.86 0.1575 0.925 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.725 0.3375 0.86 ;
        RECT 0.25 0.28 0.315 1.3725 ;
      LAYER metal2 ;
        RECT 0.27 0.725 0.34 0.86 ;
      LAYER via1 ;
        RECT 0.2725 0.76 0.3375 0.825 ;
    END
  END Y
END inv

MACRO latch
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN latch 0 0.1 ;
  SIZE 1.8925 BY 1.45 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.45 1.8925 1.65 ;
        RECT 1.5275 1.2475 1.5925 1.65 ;
        RECT 0.5925 1.22 0.6575 1.65 ;
        RECT 0.25 1.2 0.315 1.65 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 1.8925 0.2 ;
        RECT 1.5275 0 1.5925 0.385 ;
        RECT 0.5925 0 0.6575 0.385 ;
        RECT 0.25 0 0.315 0.385 ;
    END
  END vss!
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.5925 0.4525 0.6575 0.5875 ;
      LAYER metal2 ;
        RECT 0.59 0.4525 0.66 0.5875 ;
      LAYER via1 ;
        RECT 0.5925 0.4875 0.6575 0.5525 ;
    END
  END D
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.295 0.925 0.36 1.06 ;
      LAYER metal2 ;
        RECT 0.2925 0.925 0.3625 1.06 ;
      LAYER via1 ;
        RECT 0.295 0.96 0.36 1.025 ;
    END
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.7675 0.265 1.8325 1.355 ;
        RECT 1.4325 1.03 1.4975 1.165 ;
      LAYER metal2 ;
        RECT 1.765 0.89 1.835 1.355 ;
        RECT 1.4325 0.89 1.835 0.96 ;
        RECT 1.43 1.03 1.5025 1.165 ;
        RECT 1.4325 0.89 1.5025 1.165 ;
      LAYER via1 ;
        RECT 1.4325 1.065 1.4975 1.13 ;
        RECT 1.7675 1.255 1.8325 1.32 ;
    END
  END Q
  OBS
    LAYER metal1 ;
      RECT 0.78 1.22 0.845 1.355 ;
      RECT 0.7775 0.265 0.8425 1.3325 ;
      RECT 0.7775 0.265 0.845 0.4 ;
      RECT 0.06 1.2075 0.1275 1.3425 ;
      RECT 0.0625 0.265 0.1275 1.3425 ;
      RECT 0.06 0.265 0.1275 0.4 ;
      RECT 1.6275 1.03 1.6925 1.165 ;
      RECT 1.3025 0.265 1.3675 1.355 ;
      RECT 1.1725 0.405 1.2375 0.54 ;
      RECT 1.1725 0.96 1.2375 1.095 ;
      RECT 1.0425 0.265 1.1075 1.355 ;
      RECT 0.9125 0.405 0.9775 0.54 ;
      RECT 0.9125 1.015 0.9775 1.15 ;
      RECT 0.4375 0.265 0.5025 1.3425 ;
      RECT 0.195 0.47 0.26 0.605 ;
    LAYER metal2 ;
      RECT 1.04 1.43 1.69 1.5 ;
      RECT 1.62 1.03 1.69 1.5 ;
      RECT 1.04 1.22 1.11 1.5 ;
      RECT 1.62 1.03 1.695 1.165 ;
      RECT 1.17 0.96 1.24 1.095 ;
      RECT 1.1725 0.75 1.2425 1.02 ;
      RECT 1.1725 0.75 1.5 0.82 ;
      RECT 1.43 0.125 1.5 0.82 ;
      RECT 0.8825 0.405 0.98 0.54 ;
      RECT 0.8825 0.125 0.9525 0.54 ;
      RECT 0.0575 0.125 0.1275 0.4 ;
      RECT 0.0575 0.125 1.5 0.195 ;
      RECT 0.435 1.0375 0.505 1.3425 ;
      RECT 0.91 0.61 0.98 1.15 ;
      RECT 0.435 1.0375 0.98 1.1075 ;
      RECT 0.91 0.61 1.2375 0.68 ;
      RECT 1.1675 0.4275 1.2375 0.68 ;
      RECT 1.17 0.405 1.24 0.54 ;
      RECT 0.435 0.4725 0.505 0.6075 ;
      RECT 0.1925 0.47 0.2625 0.605 ;
      RECT 0.1875 0.5 0.5075 0.57 ;
    LAYER via1 ;
      RECT 1.6275 1.065 1.6925 1.13 ;
      RECT 1.1725 0.44 1.2375 0.505 ;
      RECT 1.1725 0.995 1.2375 1.06 ;
      RECT 1.0425 1.255 1.1075 1.32 ;
      RECT 0.9125 0.44 0.9775 0.505 ;
      RECT 0.9125 1.05 0.9775 1.115 ;
      RECT 0.4375 0.5075 0.5025 0.5725 ;
      RECT 0.4375 1.2425 0.5025 1.3075 ;
      RECT 0.195 0.505 0.26 0.57 ;
      RECT 0.06 0.3 0.125 0.365 ;
  END
END latch

MACRO mux2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN mux2 0 0.1 ;
  SIZE 1.6225 BY 1.45 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.45 1.6225 1.65 ;
        RECT 1.46 1.29 1.525 1.65 ;
        RECT 0.6725 1.265 0.7375 1.65 ;
        RECT 0.06 1.0225 0.125 1.65 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 1.6225 0.2 ;
        RECT 1.4975 0 1.5625 0.3625 ;
        RECT 0.6725 0 0.7375 0.415 ;
        RECT 0.06 0 0.125 0.455 ;
    END
  END vss!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.4375 0.49 1.5725 0.555 ;
        RECT 0.9625 1.0425 1.555 1.1125 ;
        RECT 1.485 0.49 1.555 1.1125 ;
        RECT 0.9325 0.9125 1.0675 0.9775 ;
        RECT 0.9625 0.9125 1.0325 1.1125 ;
      LAYER metal2 ;
        RECT 1.4375 0.4875 1.5725 0.5575 ;
      LAYER via1 ;
        RECT 1.4725 0.49 1.5375 0.555 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.72 0.9125 0.855 0.9775 ;
      LAYER metal2 ;
        RECT 0.72 0.91 0.855 0.98 ;
      LAYER via1 ;
        RECT 0.755 0.9125 0.82 0.9775 ;
    END
  END B
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.28 0.91 1.415 0.975 ;
        RECT 0.8925 0.63 1.0275 0.695 ;
        RECT 0.0375 0.735 0.1725 0.8025 ;
      LAYER metal2 ;
        RECT 1.28 0.9075 1.415 0.9775 ;
        RECT 1.3 0.6275 1.37 0.9775 ;
        RECT 0.105 0.6275 1.37 0.6975 ;
        RECT 0.0375 0.735 0.175 0.805 ;
        RECT 0.105 0.6275 0.175 0.805 ;
      LAYER via1 ;
        RECT 0.0725 0.7375 0.1375 0.8025 ;
        RECT 0.9275 0.63 0.9925 0.695 ;
        RECT 1.315 0.91 1.38 0.975 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.4175 0.275 0.4825 1.3225 ;
        RECT 0.415 0.7675 0.4825 0.9025 ;
      LAYER metal2 ;
        RECT 0.4125 0.7675 0.4825 0.9025 ;
      LAYER via1 ;
        RECT 0.415 0.8025 0.48 0.8675 ;
    END
  END Y
  OBS
    LAYER metal1 ;
      RECT 0.9725 0.7725 1.1625 0.8375 ;
      RECT 1.0975 0.3125 1.1625 0.8375 ;
      RECT 0.975 0.77 1.1625 0.8375 ;
      RECT 1.05 0.2775 1.115 0.4125 ;
      RECT 0.25 0.29 0.315 1.355 ;
      RECT 0.21 0.49 0.345 0.555 ;
      RECT 1.2325 0.49 1.3675 0.555 ;
      RECT 1.27 1.185 1.335 1.32 ;
      RECT 1.0475 1.18 1.1825 1.245 ;
      RECT 0.86 1.185 0.925 1.32 ;
      RECT 0.5525 0.77 0.6875 0.835 ;
    LAYER metal2 ;
      RECT 0.8575 1.3175 1.3375 1.3875 ;
      RECT 1.2675 1.185 1.3375 1.3875 ;
      RECT 0.8575 1.185 0.9275 1.3875 ;
      RECT 1.0475 1.1775 1.1825 1.2475 ;
      RECT 1.08 0.7675 1.15 1.2475 ;
      RECT 0.5525 0.7675 1.15 0.8375 ;
      RECT 0.1825 0.4875 1.3675 0.5575 ;
    LAYER via1 ;
      RECT 1.27 1.22 1.335 1.285 ;
      RECT 1.2675 0.49 1.3325 0.555 ;
      RECT 1.0825 1.18 1.1475 1.245 ;
      RECT 1.01 0.77 1.075 0.835 ;
      RECT 0.86 1.22 0.925 1.285 ;
      RECT 0.5875 0.77 0.6525 0.835 ;
      RECT 0.245 0.49 0.31 0.555 ;
  END
END mux2

MACRO nand2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN nand2 0 0.1 ;
  SIZE 0.56 BY 1.45 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.45 0.56 1.65 ;
        RECT 0.435 1.0575 0.5 1.65 ;
        RECT 0.06 1.0375 0.125 1.65 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.56 0.2 ;
        RECT 0.06 0 0.125 0.4225 ;
    END
  END vss!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.05 0.79 0.185 0.855 ;
      LAYER metal2 ;
        RECT 0.05 0.7875 0.185 0.8575 ;
      LAYER via1 ;
        RECT 0.085 0.79 0.15 0.855 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.255 0.785 0.39 0.85 ;
      LAYER metal2 ;
        RECT 0.255 0.7825 0.39 0.8525 ;
      LAYER via1 ;
        RECT 0.29 0.785 0.355 0.85 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2475 0.915 0.52 0.98 ;
        RECT 0.455 0.28 0.52 0.98 ;
        RECT 0.435 0.2775 0.5 0.485 ;
        RECT 0.2475 0.915 0.3125 1.155 ;
      LAYER metal2 ;
        RECT 0.245 0.925 0.315 1.06 ;
      LAYER via1 ;
        RECT 0.2475 0.96 0.3125 1.025 ;
    END
  END Y
END nand2

MACRO nor2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN nor2 0 0.1 ;
  SIZE 0.56 BY 1.45 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.45 0.56 1.65 ;
        RECT 0.06 1.0375 0.125 1.65 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.56 0.2 ;
        RECT 0.435 0 0.5 0.385 ;
        RECT 0.06 0 0.125 0.3975 ;
    END
  END vss!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.035 0.9075 0.17 0.9725 ;
      LAYER metal2 ;
        RECT 0.035 0.905 0.17 0.975 ;
      LAYER via1 ;
        RECT 0.07 0.9075 0.135 0.9725 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.39 0.545 0.455 0.68 ;
      LAYER metal2 ;
        RECT 0.3875 0.545 0.4575 0.68 ;
      LAYER via1 ;
        RECT 0.39 0.58 0.455 0.645 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.455 0.8 0.5225 0.935 ;
        RECT 0.435 1.0575 0.52 1.1925 ;
        RECT 0.455 0.7775 0.52 1.1925 ;
        RECT 0.2475 0.7775 0.52 0.8425 ;
        RECT 0.2475 0.265 0.3125 0.8425 ;
      LAYER metal2 ;
        RECT 0.455 0.8 0.525 0.935 ;
      LAYER via1 ;
        RECT 0.4575 0.835 0.5225 0.9 ;
    END
  END Y
END nor2

MACRO oai21
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN oai21 0 0.1 ;
  SIZE 0.75 BY 1.45 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.45 0.75 1.65 ;
        RECT 0.625 1.2525 0.69 1.65 ;
        RECT 0.06 1.065 0.125 1.65 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.75 0.2 ;
        RECT 0.06 0 0.125 0.4125 ;
    END
  END vss!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.5 0.7325 0.565 0.8675 ;
      LAYER metal2 ;
        RECT 0.4975 0.7325 0.5675 0.8675 ;
      LAYER via1 ;
        RECT 0.5 0.7675 0.565 0.8325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.3075 0.7375 0.3725 0.8725 ;
      LAYER metal2 ;
        RECT 0.305 0.7375 0.375 0.8725 ;
      LAYER via1 ;
        RECT 0.3075 0.7725 0.3725 0.8375 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.1025 0.7375 0.1675 0.8725 ;
      LAYER metal2 ;
        RECT 0.1 0.7375 0.17 0.8725 ;
      LAYER via1 ;
        RECT 0.1025 0.7725 0.1675 0.8375 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2475 0.995 0.715 1.06 ;
        RECT 0.65 0.5175 0.715 1.06 ;
        RECT 0.6475 0.7375 0.715 0.8725 ;
        RECT 0.4375 0.5175 0.715 0.5825 ;
        RECT 0.4375 0.265 0.5025 0.5825 ;
        RECT 0.2475 0.995 0.3125 1.2075 ;
      LAYER metal2 ;
        RECT 0.645 0.7375 0.715 0.8725 ;
        RECT 0.245 1.0725 0.315 1.2075 ;
      LAYER via1 ;
        RECT 0.2475 1.1075 0.3125 1.1725 ;
        RECT 0.6475 0.7725 0.7125 0.8375 ;
    END
  END Y
  OBS
    LAYER metal1 ;
      RECT 0.625 0.265 0.69 0.4 ;
      RECT 0.2475 0.265 0.3125 0.4125 ;
    LAYER metal2 ;
      RECT 0.245 0.435 0.6925 0.505 ;
      RECT 0.6225 0.265 0.6925 0.505 ;
      RECT 0.245 0.26 0.315 0.505 ;
    LAYER via1 ;
      RECT 0.625 0.3 0.69 0.365 ;
      RECT 0.2475 0.3075 0.3125 0.3725 ;
  END
END oai21

MACRO or2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN or2 0 0.1 ;
  SIZE 0.8 BY 1.45 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.45 0.8 1.65 ;
        RECT 0.3 1.2175 0.365 1.65 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 0.8 0.2 ;
        RECT 0.675 0 0.74 0.385 ;
        RECT 0.3 0 0.365 0.385 ;
    END
  END vss!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.29 0.915 0.425 0.98 ;
      LAYER metal2 ;
        RECT 0.29 0.9125 0.425 0.9825 ;
      LAYER via1 ;
        RECT 0.325 0.915 0.39 0.98 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.495 0.9125 0.63 0.9775 ;
      LAYER metal2 ;
        RECT 0.495 0.91 0.63 0.98 ;
      LAYER via1 ;
        RECT 0.53 0.9125 0.595 0.9775 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.265 0.125 1.2325 ;
        RECT 0.0375 0.785 0.125 0.92 ;
      LAYER metal2 ;
        RECT 0.035 0.785 0.105 0.92 ;
      LAYER via1 ;
        RECT 0.0375 0.82 0.1025 0.885 ;
    END
  END Y
  OBS
    LAYER metal1 ;
      RECT 0.675 1.1225 0.765 1.2575 ;
      RECT 0.7 0.7775 0.765 1.2575 ;
      RECT 0.4875 0.7775 0.765 0.8425 ;
      RECT 0.1925 0.765 0.5525 0.83 ;
      RECT 0.4875 0.265 0.5525 0.8425 ;
  END
END or2

MACRO xnor2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN xnor2 0 0.1 ;
  SIZE 1.205 BY 1.45 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.45 1.205 1.65 ;
        RECT 1.08 1.29 1.145 1.65 ;
        RECT 0.515 1.2175 0.58 1.65 ;
        RECT 0.095 1.27 0.16 1.65 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 1.205 0.2 ;
        RECT 0.515 0 0.58 0.36 ;
    END
  END vss!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.955 0.83 1.02 0.965 ;
        RECT 0.4225 1.025 1.0075 1.09 ;
        RECT 0.9425 0.86 1.0075 1.09 ;
        RECT 0.4225 0.8225 0.4875 1.09 ;
        RECT 0.42 0.8175 0.485 0.9525 ;
      LAYER metal2 ;
        RECT 0.9525 0.83 1.0225 0.965 ;
        RECT 0.4175 0.8175 0.4875 0.9525 ;
      LAYER via1 ;
        RECT 0.42 0.8525 0.485 0.9175 ;
        RECT 0.955 0.865 1.02 0.93 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.745 0.8175 0.81 0.9525 ;
        RECT 0.0775 0.89 0.2125 0.955 ;
      LAYER metal2 ;
        RECT 0.1425 1.0225 0.8175 1.0925 ;
        RECT 0.7475 0.865 0.8175 1.0925 ;
        RECT 0.7425 0.8175 0.8125 0.9525 ;
        RECT 0.1425 0.885 0.2125 1.0925 ;
        RECT 0.0775 0.8875 0.2125 0.9575 ;
      LAYER via1 ;
        RECT 0.1125 0.89 0.1775 0.955 ;
        RECT 0.745 0.8525 0.81 0.9175 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.7025 1.16 1.17 1.225 ;
        RECT 1.105 0.6375 1.17 1.225 ;
        RECT 1.1025 0.8375 1.17 0.9725 ;
        RECT 0.8925 0.6375 1.17 0.7025 ;
        RECT 0.8925 0.265 0.9575 0.7025 ;
        RECT 0.7025 1.16 0.7675 1.36 ;
      LAYER metal2 ;
        RECT 1.1 0.8375 1.17 0.9725 ;
        RECT 0.7 1.225 0.77 1.36 ;
      LAYER via1 ;
        RECT 0.7025 1.26 0.7675 1.325 ;
        RECT 1.1025 0.8725 1.1675 0.9375 ;
    END
  END Y
  OBS
    LAYER metal1 ;
      RECT 0.2825 0.6875 0.3475 1.385 ;
      RECT 0.57 0.6875 0.635 0.95 ;
      RECT 0.095 0.6875 0.635 0.7525 ;
      RECT 0.095 0.265 0.16 0.7525 ;
      RECT 1.08 0.265 1.145 0.4 ;
      RECT 0.7025 0.265 0.7675 0.4125 ;
    LAYER metal2 ;
      RECT 0.7 0.2 0.77 0.4125 ;
      RECT 1.075 0.265 1.1475 0.4 ;
      RECT 0.7 0.2 1.145 0.27 ;
    LAYER via1 ;
      RECT 1.08 0.3 1.145 0.365 ;
      RECT 0.7025 0.3075 0.7675 0.3725 ;
  END
END xnor2

MACRO xor2
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN xor2 0 0.1 ;
  SIZE 1.28 BY 1.45 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.45 1.28 1.65 ;
        RECT 0.59 1.2675 0.655 1.65 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 0 1.28 0.2 ;
        RECT 1.155 0 1.22 0.36 ;
        RECT 0.59 0 0.655 0.385 ;
        RECT 0.06 0 0.125 0.3975 ;
    END
  END vss!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.19 1.04 0.9025 1.105 ;
        RECT 0.8375 0.895 0.9025 1.105 ;
        RECT 0.82 0.8125 0.885 0.9475 ;
        RECT 0.19 0.8175 0.255 1.105 ;
        RECT 0.1825 0.8125 0.2475 0.9475 ;
      LAYER metal2 ;
        RECT 0.8175 0.8125 0.8875 0.9475 ;
        RECT 0.18 0.8125 0.25 0.9475 ;
      LAYER via1 ;
        RECT 0.1825 0.8475 0.2475 0.9125 ;
        RECT 0.82 0.8475 0.885 0.9125 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.03 0.8125 1.095 0.9475 ;
        RECT 0.3875 0.8125 0.4525 0.9475 ;
      LAYER metal2 ;
        RECT 1.0275 0.8125 1.0975 0.9475 ;
        RECT 0.995 0.48 1.065 0.9275 ;
        RECT 0.3875 0.48 1.065 0.55 ;
        RECT 0.3875 0.48 0.4575 0.9125 ;
        RECT 0.385 0.8125 0.455 0.9475 ;
      LAYER via1 ;
        RECT 0.3875 0.8475 0.4525 0.9125 ;
        RECT 1.03 0.8475 1.095 0.9125 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.9675 1.04 1.245 1.105 ;
        RECT 1.18 0.4725 1.245 1.105 ;
        RECT 1.175 0.79 1.245 0.925 ;
        RECT 0.7775 0.4725 1.245 0.5375 ;
        RECT 0.9675 1.04 1.0325 1.2175 ;
        RECT 0.7775 0.265 0.8425 0.5375 ;
      LAYER metal2 ;
        RECT 1.1725 0.79 1.2425 0.925 ;
      LAYER via1 ;
        RECT 1.175 0.825 1.24 0.89 ;
    END
  END Y
  OBS
    LAYER metal1 ;
      RECT 0.035 0.5375 0.1 1.195 ;
      RECT 0.035 1.0575 0.125 1.1925 ;
      RECT 0.6375 0.8125 0.7025 0.9475 ;
      RECT 0.5925 0.5375 0.6575 0.925 ;
      RECT 0.035 0.5375 0.6575 0.6025 ;
      RECT 0.2475 0.265 0.3125 0.6025 ;
      RECT 1.155 1.1725 1.22 1.3125 ;
      RECT 0.7775 1.18 0.8425 1.32 ;
    LAYER metal2 ;
      RECT 0.7725 1.2975 1.2225 1.3675 ;
      RECT 1.1525 1.1725 1.2225 1.3675 ;
      RECT 0.7725 1.185 0.845 1.3675 ;
      RECT 0.7725 1.18 0.8425 1.3675 ;
      RECT 0.635 0.8125 0.705 0.9475 ;
    LAYER via1 ;
      RECT 1.155 1.2125 1.22 1.2775 ;
      RECT 0.7775 1.22 0.8425 1.285 ;
      RECT 0.6375 0.8475 0.7025 0.9125 ;
  END
END xor2

END LIBRARY
