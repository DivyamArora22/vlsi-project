VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO regfile
  CLASS CORE ;
  ORIGIN 0 -0.1 ;
  FOREIGN regfile 0 0.1 ;
  SIZE 115.435 BY 1.45 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.45 115.435 1.65 ;
        RECT 115.07 1.2475 115.135 1.65 ;
        RECT 114.135 1.22 114.2 1.65 ;
        RECT 113.7925 1.2 113.8575 1.65 ;
        RECT 113.2275 1.2 113.2925 1.65 ;
        RECT 112.885 1.22 112.95 1.65 ;
        RECT 111.95 1.2475 112.015 1.65 ;
        RECT 111.325 1.23 111.39 1.65 ;
        RECT 110.94 1.23 111.005 1.65 ;
        RECT 110.755 1.05 110.82 1.65 ;
        RECT 110.37 1.05 110.435 1.65 ;
        RECT 109.215 1.23 109.28 1.65 ;
        RECT 108.63 1.23 108.695 1.65 ;
        RECT 107.475 1.05 107.54 1.65 ;
        RECT 107.29 1.05 107.355 1.65 ;
        RECT 106.905 1.05 106.97 1.65 ;
        RECT 105.75 1.23 105.815 1.65 ;
        RECT 105.165 1.23 105.23 1.65 ;
        RECT 104.01 1.05 104.075 1.65 ;
        RECT 103.825 1.05 103.89 1.65 ;
        RECT 103.44 1.05 103.505 1.65 ;
        RECT 102.285 1.23 102.35 1.65 ;
        RECT 101.7 1.23 101.765 1.65 ;
        RECT 100.545 1.05 100.61 1.65 ;
        RECT 100.36 1.05 100.425 1.65 ;
        RECT 99.975 1.05 100.04 1.65 ;
        RECT 98.82 1.23 98.885 1.65 ;
        RECT 98.235 1.23 98.3 1.65 ;
        RECT 97.08 1.05 97.145 1.65 ;
        RECT 96.895 1.05 96.96 1.65 ;
        RECT 96.51 1.05 96.575 1.65 ;
        RECT 95.355 1.23 95.42 1.65 ;
        RECT 94.77 1.23 94.835 1.65 ;
        RECT 93.615 1.05 93.68 1.65 ;
        RECT 93.43 1.05 93.495 1.65 ;
        RECT 93.045 1.05 93.11 1.65 ;
        RECT 91.89 1.23 91.955 1.65 ;
        RECT 91.305 1.23 91.37 1.65 ;
        RECT 90.15 1.05 90.215 1.65 ;
        RECT 89.965 1.05 90.03 1.65 ;
        RECT 89.58 1.05 89.645 1.65 ;
        RECT 88.425 1.23 88.49 1.65 ;
        RECT 87.84 1.23 87.905 1.65 ;
        RECT 86.685 1.05 86.75 1.65 ;
        RECT 86.5 1.05 86.565 1.65 ;
        RECT 86.115 1.05 86.18 1.65 ;
        RECT 84.96 1.23 85.025 1.65 ;
        RECT 84.375 1.23 84.44 1.65 ;
        RECT 83.22 1.05 83.285 1.65 ;
        RECT 83.035 1.05 83.1 1.65 ;
        RECT 82.65 1.05 82.715 1.65 ;
        RECT 81.495 1.23 81.56 1.65 ;
        RECT 80.91 1.23 80.975 1.65 ;
        RECT 79.755 1.05 79.82 1.65 ;
        RECT 79.57 1.05 79.635 1.65 ;
        RECT 79.185 1.05 79.25 1.65 ;
        RECT 78.03 1.23 78.095 1.65 ;
        RECT 77.445 1.23 77.51 1.65 ;
        RECT 76.29 1.05 76.355 1.65 ;
        RECT 76.105 1.05 76.17 1.65 ;
        RECT 75.72 1.05 75.785 1.65 ;
        RECT 74.565 1.23 74.63 1.65 ;
        RECT 73.98 1.23 74.045 1.65 ;
        RECT 72.825 1.05 72.89 1.65 ;
        RECT 72.64 1.05 72.705 1.65 ;
        RECT 72.255 1.05 72.32 1.65 ;
        RECT 71.1 1.23 71.165 1.65 ;
        RECT 70.515 1.23 70.58 1.65 ;
        RECT 69.36 1.05 69.425 1.65 ;
        RECT 69.175 1.05 69.24 1.65 ;
        RECT 68.79 1.05 68.855 1.65 ;
        RECT 67.635 1.23 67.7 1.65 ;
        RECT 67.05 1.23 67.115 1.65 ;
        RECT 65.895 1.05 65.96 1.65 ;
        RECT 65.71 1.05 65.775 1.65 ;
        RECT 65.325 1.05 65.39 1.65 ;
        RECT 64.17 1.23 64.235 1.65 ;
        RECT 63.585 1.23 63.65 1.65 ;
        RECT 62.43 1.05 62.495 1.65 ;
        RECT 62.245 1.05 62.31 1.65 ;
        RECT 61.86 1.05 61.925 1.65 ;
        RECT 60.705 1.23 60.77 1.65 ;
        RECT 60.12 1.23 60.185 1.65 ;
        RECT 58.965 1.05 59.03 1.65 ;
        RECT 58.78 1.05 58.845 1.65 ;
        RECT 58.395 1.05 58.46 1.65 ;
        RECT 57.24 1.23 57.305 1.65 ;
        RECT 56.655 1.23 56.72 1.65 ;
        RECT 55.5 1.05 55.565 1.65 ;
        RECT 55.315 1.05 55.38 1.65 ;
        RECT 54.93 1.05 54.995 1.65 ;
        RECT 53.775 1.23 53.84 1.65 ;
        RECT 53.19 1.23 53.255 1.65 ;
        RECT 52.035 1.05 52.1 1.65 ;
        RECT 51.85 1.05 51.915 1.65 ;
        RECT 51.465 1.05 51.53 1.65 ;
        RECT 50.31 1.23 50.375 1.65 ;
        RECT 49.725 1.23 49.79 1.65 ;
        RECT 48.57 1.05 48.635 1.65 ;
        RECT 48.385 1.05 48.45 1.65 ;
        RECT 48 1.05 48.065 1.65 ;
        RECT 46.845 1.23 46.91 1.65 ;
        RECT 46.26 1.23 46.325 1.65 ;
        RECT 45.105 1.05 45.17 1.65 ;
        RECT 44.92 1.05 44.985 1.65 ;
        RECT 44.535 1.05 44.6 1.65 ;
        RECT 43.38 1.23 43.445 1.65 ;
        RECT 42.795 1.23 42.86 1.65 ;
        RECT 41.64 1.05 41.705 1.65 ;
        RECT 41.455 1.05 41.52 1.65 ;
        RECT 41.07 1.05 41.135 1.65 ;
        RECT 39.915 1.23 39.98 1.65 ;
        RECT 39.33 1.23 39.395 1.65 ;
        RECT 38.175 1.05 38.24 1.65 ;
        RECT 37.99 1.05 38.055 1.65 ;
        RECT 37.605 1.05 37.67 1.65 ;
        RECT 36.45 1.23 36.515 1.65 ;
        RECT 35.865 1.23 35.93 1.65 ;
        RECT 34.71 1.05 34.775 1.65 ;
        RECT 34.525 1.05 34.59 1.65 ;
        RECT 34.14 1.05 34.205 1.65 ;
        RECT 32.985 1.23 33.05 1.65 ;
        RECT 32.4 1.23 32.465 1.65 ;
        RECT 31.245 1.05 31.31 1.65 ;
        RECT 31.06 1.05 31.125 1.65 ;
        RECT 30.675 1.05 30.74 1.65 ;
        RECT 29.52 1.23 29.585 1.65 ;
        RECT 28.935 1.23 29 1.65 ;
        RECT 27.78 1.05 27.845 1.65 ;
        RECT 27.595 1.05 27.66 1.65 ;
        RECT 27.21 1.05 27.275 1.65 ;
        RECT 26.055 1.23 26.12 1.65 ;
        RECT 25.47 1.23 25.535 1.65 ;
        RECT 24.315 1.05 24.38 1.65 ;
        RECT 24.13 1.05 24.195 1.65 ;
        RECT 23.745 1.05 23.81 1.65 ;
        RECT 22.59 1.23 22.655 1.65 ;
        RECT 22.005 1.23 22.07 1.65 ;
        RECT 20.85 1.05 20.915 1.65 ;
        RECT 20.665 1.05 20.73 1.65 ;
        RECT 20.28 1.05 20.345 1.65 ;
        RECT 19.125 1.23 19.19 1.65 ;
        RECT 18.54 1.23 18.605 1.65 ;
        RECT 17.385 1.05 17.45 1.65 ;
        RECT 17.2 1.05 17.265 1.65 ;
        RECT 16.815 1.05 16.88 1.65 ;
        RECT 15.66 1.23 15.725 1.65 ;
        RECT 15.075 1.23 15.14 1.65 ;
        RECT 13.92 1.05 13.985 1.65 ;
        RECT 13.735 1.05 13.8 1.65 ;
        RECT 13.35 1.05 13.415 1.65 ;
        RECT 12.195 1.23 12.26 1.65 ;
        RECT 11.61 1.23 11.675 1.65 ;
        RECT 10.455 1.05 10.52 1.65 ;
        RECT 10.27 1.05 10.335 1.65 ;
        RECT 9.885 1.05 9.95 1.65 ;
        RECT 8.73 1.23 8.795 1.65 ;
        RECT 8.145 1.23 8.21 1.65 ;
        RECT 6.99 1.05 7.055 1.65 ;
        RECT 6.805 1.05 6.87 1.65 ;
        RECT 6.42 1.05 6.485 1.65 ;
        RECT 5.265 1.23 5.33 1.65 ;
        RECT 4.68 1.23 4.745 1.65 ;
        RECT 3.525 1.05 3.59 1.65 ;
        RECT 3.34 1.05 3.405 1.65 ;
        RECT 2.955 1.05 3.02 1.65 ;
        RECT 1.8 1.23 1.865 1.65 ;
        RECT 1.215 1.23 1.28 1.65 ;
        RECT 0.06 1.05 0.125 1.65 ;
    END
  END vdd!
  PIN vss!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
        RECT 0.425 0.845 0.495 0.985 ;
      LAYER metal1 ;
        RECT 0 0 115.435 0.2 ;
        RECT 115.07 0 115.135 0.385 ;
        RECT 114.135 0 114.2 0.385 ;
        RECT 113.7925 0 113.8575 0.385 ;
        RECT 113.2275 0 113.2925 0.385 ;
        RECT 112.885 0 112.95 0.385 ;
        RECT 111.95 0 112.015 0.385 ;
        RECT 111.325 0 111.39 0.39 ;
        RECT 110.94 0 111.005 0.415 ;
        RECT 110.755 0 110.82 0.39 ;
        RECT 110.37 0 110.435 0.415 ;
        RECT 109.215 0 109.28 0.415 ;
        RECT 108.63 0 108.695 0.415 ;
        RECT 107.475 0 107.54 0.415 ;
        RECT 107.29 0 107.355 0.39 ;
        RECT 106.905 0 106.97 0.415 ;
        RECT 105.75 0 105.815 0.415 ;
        RECT 105.165 0 105.23 0.415 ;
        RECT 104.01 0 104.075 0.415 ;
        RECT 103.825 0 103.89 0.39 ;
        RECT 103.44 0 103.505 0.415 ;
        RECT 102.285 0 102.35 0.415 ;
        RECT 101.7 0 101.765 0.415 ;
        RECT 100.545 0 100.61 0.415 ;
        RECT 100.36 0 100.425 0.39 ;
        RECT 99.975 0 100.04 0.415 ;
        RECT 98.82 0 98.885 0.415 ;
        RECT 98.235 0 98.3 0.415 ;
        RECT 97.08 0 97.145 0.415 ;
        RECT 96.895 0 96.96 0.39 ;
        RECT 96.51 0 96.575 0.415 ;
        RECT 95.355 0 95.42 0.415 ;
        RECT 94.77 0 94.835 0.415 ;
        RECT 93.615 0 93.68 0.415 ;
        RECT 93.43 0 93.495 0.39 ;
        RECT 93.045 0 93.11 0.415 ;
        RECT 91.89 0 91.955 0.415 ;
        RECT 91.305 0 91.37 0.415 ;
        RECT 90.15 0 90.215 0.415 ;
        RECT 89.965 0 90.03 0.39 ;
        RECT 89.58 0 89.645 0.415 ;
        RECT 88.425 0 88.49 0.415 ;
        RECT 87.84 0 87.905 0.415 ;
        RECT 86.685 0 86.75 0.415 ;
        RECT 86.5 0 86.565 0.39 ;
        RECT 86.115 0 86.18 0.415 ;
        RECT 84.96 0 85.025 0.415 ;
        RECT 84.375 0 84.44 0.415 ;
        RECT 83.22 0 83.285 0.415 ;
        RECT 83.035 0 83.1 0.39 ;
        RECT 82.65 0 82.715 0.415 ;
        RECT 81.495 0 81.56 0.415 ;
        RECT 80.91 0 80.975 0.415 ;
        RECT 79.755 0 79.82 0.415 ;
        RECT 79.57 0 79.635 0.39 ;
        RECT 79.185 0 79.25 0.415 ;
        RECT 78.03 0 78.095 0.415 ;
        RECT 77.445 0 77.51 0.415 ;
        RECT 76.29 0 76.355 0.415 ;
        RECT 76.105 0 76.17 0.39 ;
        RECT 75.72 0 75.785 0.415 ;
        RECT 74.565 0 74.63 0.415 ;
        RECT 73.98 0 74.045 0.415 ;
        RECT 72.825 0 72.89 0.415 ;
        RECT 72.64 0 72.705 0.39 ;
        RECT 72.255 0 72.32 0.415 ;
        RECT 71.1 0 71.165 0.415 ;
        RECT 70.515 0 70.58 0.415 ;
        RECT 69.36 0 69.425 0.415 ;
        RECT 69.175 0 69.24 0.39 ;
        RECT 68.79 0 68.855 0.415 ;
        RECT 67.635 0 67.7 0.415 ;
        RECT 67.05 0 67.115 0.415 ;
        RECT 65.895 0 65.96 0.415 ;
        RECT 65.71 0 65.775 0.39 ;
        RECT 65.325 0 65.39 0.415 ;
        RECT 64.17 0 64.235 0.415 ;
        RECT 63.585 0 63.65 0.415 ;
        RECT 62.43 0 62.495 0.415 ;
        RECT 62.245 0 62.31 0.39 ;
        RECT 61.86 0 61.925 0.415 ;
        RECT 60.705 0 60.77 0.415 ;
        RECT 60.12 0 60.185 0.415 ;
        RECT 58.965 0 59.03 0.415 ;
        RECT 58.78 0 58.845 0.39 ;
        RECT 58.395 0 58.46 0.415 ;
        RECT 57.24 0 57.305 0.415 ;
        RECT 56.655 0 56.72 0.415 ;
        RECT 55.5 0 55.565 0.415 ;
        RECT 55.315 0 55.38 0.39 ;
        RECT 54.93 0 54.995 0.415 ;
        RECT 53.775 0 53.84 0.415 ;
        RECT 53.19 0 53.255 0.415 ;
        RECT 52.035 0 52.1 0.415 ;
        RECT 51.85 0 51.915 0.39 ;
        RECT 51.465 0 51.53 0.415 ;
        RECT 50.31 0 50.375 0.415 ;
        RECT 49.725 0 49.79 0.415 ;
        RECT 48.57 0 48.635 0.415 ;
        RECT 48.385 0 48.45 0.39 ;
        RECT 48 0 48.065 0.415 ;
        RECT 46.845 0 46.91 0.415 ;
        RECT 46.26 0 46.325 0.415 ;
        RECT 45.105 0 45.17 0.415 ;
        RECT 44.92 0 44.985 0.39 ;
        RECT 44.535 0 44.6 0.415 ;
        RECT 43.38 0 43.445 0.415 ;
        RECT 42.795 0 42.86 0.415 ;
        RECT 41.64 0 41.705 0.415 ;
        RECT 41.455 0 41.52 0.39 ;
        RECT 41.07 0 41.135 0.415 ;
        RECT 39.915 0 39.98 0.415 ;
        RECT 39.33 0 39.395 0.415 ;
        RECT 38.175 0 38.24 0.415 ;
        RECT 37.99 0 38.055 0.39 ;
        RECT 37.605 0 37.67 0.415 ;
        RECT 36.45 0 36.515 0.415 ;
        RECT 35.865 0 35.93 0.415 ;
        RECT 34.71 0 34.775 0.415 ;
        RECT 34.525 0 34.59 0.39 ;
        RECT 34.14 0 34.205 0.415 ;
        RECT 32.985 0 33.05 0.415 ;
        RECT 32.4 0 32.465 0.415 ;
        RECT 31.245 0 31.31 0.415 ;
        RECT 31.06 0 31.125 0.39 ;
        RECT 30.675 0 30.74 0.415 ;
        RECT 29.52 0 29.585 0.415 ;
        RECT 28.935 0 29 0.415 ;
        RECT 27.78 0 27.845 0.415 ;
        RECT 27.595 0 27.66 0.39 ;
        RECT 27.21 0 27.275 0.415 ;
        RECT 26.055 0 26.12 0.415 ;
        RECT 25.47 0 25.535 0.415 ;
        RECT 24.315 0 24.38 0.415 ;
        RECT 24.13 0 24.195 0.39 ;
        RECT 23.745 0 23.81 0.415 ;
        RECT 22.59 0 22.655 0.415 ;
        RECT 22.005 0 22.07 0.415 ;
        RECT 20.85 0 20.915 0.415 ;
        RECT 20.665 0 20.73 0.39 ;
        RECT 20.28 0 20.345 0.415 ;
        RECT 19.125 0 19.19 0.415 ;
        RECT 18.54 0 18.605 0.415 ;
        RECT 17.385 0 17.45 0.415 ;
        RECT 17.2 0 17.265 0.39 ;
        RECT 16.815 0 16.88 0.415 ;
        RECT 15.66 0 15.725 0.415 ;
        RECT 15.075 0 15.14 0.415 ;
        RECT 13.92 0 13.985 0.415 ;
        RECT 13.735 0 13.8 0.39 ;
        RECT 13.35 0 13.415 0.415 ;
        RECT 12.195 0 12.26 0.415 ;
        RECT 11.61 0 11.675 0.415 ;
        RECT 10.455 0 10.52 0.415 ;
        RECT 10.27 0 10.335 0.39 ;
        RECT 9.885 0 9.95 0.415 ;
        RECT 8.73 0 8.795 0.415 ;
        RECT 8.145 0 8.21 0.415 ;
        RECT 6.99 0 7.055 0.415 ;
        RECT 6.805 0 6.87 0.39 ;
        RECT 6.42 0 6.485 0.415 ;
        RECT 5.265 0 5.33 0.415 ;
        RECT 4.68 0 4.745 0.415 ;
        RECT 3.525 0 3.59 0.415 ;
        RECT 3.34 0 3.405 0.39 ;
        RECT 2.955 0 3.02 0.415 ;
        RECT 1.8 0 1.865 0.415 ;
        RECT 1.215 0 1.28 0.415 ;
        RECT 0.445 0.4875 0.51 1.14 ;
        RECT 0.4125 0 0.4775 0.985 ;
        RECT 0.06 0 0.125 0.415 ;
      LAYER metal2 ;
        RECT 0.425 0.845 0.495 0.985 ;
      LAYER via2 ;
        RECT 0.425 0.88 0.495 0.95 ;
      LAYER via1 ;
        RECT 0.4275 0.8825 0.4925 0.9475 ;
    END
  END vss!
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 113.8375 0.925 113.9025 1.06 ;
        RECT 113.1825 0.925 113.2475 1.06 ;
      LAYER metal2 ;
        RECT 113.835 0.925 113.905 1.06 ;
        RECT 113.18 0.9575 113.905 1.0275 ;
        RECT 113.18 0.925 113.25 1.06 ;
      LAYER via1 ;
        RECT 113.1825 0.96 113.2475 1.025 ;
        RECT 113.8375 0.96 113.9025 1.025 ;
    END
  END clk
  PIN rd_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.1175 0.82 0.1875 0.96 ;
      LAYER metal1 ;
        RECT 0.9025 1.2725 1.0375 1.3375 ;
        RECT 0.5425 0.2825 0.6075 0.4175 ;
        RECT 0.12 0.825 0.185 0.96 ;
      LAYER metal2 ;
        RECT 0.9025 1.27 1.0375 1.34 ;
        RECT 0.1175 1.455 0.995 1.525 ;
        RECT 0.925 1.2675 0.995 1.525 ;
        RECT 0.1175 0.4025 0.61 0.4725 ;
        RECT 0.54 0.2825 0.61 0.4725 ;
        RECT 0.1175 0.4025 0.1875 1.525 ;
      LAYER via1 ;
        RECT 0.12 0.86 0.185 0.925 ;
        RECT 0.5425 0.3175 0.6075 0.3825 ;
        RECT 0.9375 1.2725 1.0025 1.3375 ;
      LAYER via2 ;
        RECT 0.1175 0.855 0.1875 0.925 ;
    END
  END rd_sel[0]
  PIN rd_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 34.7675 0.82 34.8375 0.96 ;
      LAYER metal1 ;
        RECT 35.5525 1.2725 35.6875 1.3375 ;
        RECT 35.1925 0.2825 35.2575 0.4175 ;
        RECT 34.77 0.825 34.835 0.96 ;
      LAYER metal2 ;
        RECT 35.5525 1.27 35.6875 1.34 ;
        RECT 34.7675 1.455 35.645 1.525 ;
        RECT 35.575 1.2675 35.645 1.525 ;
        RECT 34.7675 0.4025 35.26 0.4725 ;
        RECT 35.19 0.2825 35.26 0.4725 ;
        RECT 34.7675 0.4025 34.8375 1.525 ;
      LAYER via1 ;
        RECT 34.77 0.86 34.835 0.925 ;
        RECT 35.1925 0.3175 35.2575 0.3825 ;
        RECT 35.5875 1.2725 35.6525 1.3375 ;
      LAYER via2 ;
        RECT 34.7675 0.855 34.8375 0.925 ;
    END
  END rd_sel[10]
  PIN rd_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 38.2325 0.82 38.3025 0.96 ;
      LAYER metal1 ;
        RECT 39.0175 1.2725 39.1525 1.3375 ;
        RECT 38.6575 0.2825 38.7225 0.4175 ;
        RECT 38.235 0.825 38.3 0.96 ;
      LAYER metal2 ;
        RECT 39.0175 1.27 39.1525 1.34 ;
        RECT 38.2325 1.455 39.11 1.525 ;
        RECT 39.04 1.2675 39.11 1.525 ;
        RECT 38.2325 0.4025 38.725 0.4725 ;
        RECT 38.655 0.2825 38.725 0.4725 ;
        RECT 38.2325 0.4025 38.3025 1.525 ;
      LAYER via1 ;
        RECT 38.235 0.86 38.3 0.925 ;
        RECT 38.6575 0.3175 38.7225 0.3825 ;
        RECT 39.0525 1.2725 39.1175 1.3375 ;
      LAYER via2 ;
        RECT 38.2325 0.855 38.3025 0.925 ;
    END
  END rd_sel[11]
  PIN rd_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 41.6975 0.82 41.7675 0.96 ;
      LAYER metal1 ;
        RECT 42.4825 1.2725 42.6175 1.3375 ;
        RECT 42.1225 0.2825 42.1875 0.4175 ;
        RECT 41.7 0.825 41.765 0.96 ;
      LAYER metal2 ;
        RECT 42.4825 1.27 42.6175 1.34 ;
        RECT 41.6975 1.455 42.575 1.525 ;
        RECT 42.505 1.2675 42.575 1.525 ;
        RECT 41.6975 0.4025 42.19 0.4725 ;
        RECT 42.12 0.2825 42.19 0.4725 ;
        RECT 41.6975 0.4025 41.7675 1.525 ;
      LAYER via1 ;
        RECT 41.7 0.86 41.765 0.925 ;
        RECT 42.1225 0.3175 42.1875 0.3825 ;
        RECT 42.5175 1.2725 42.5825 1.3375 ;
      LAYER via2 ;
        RECT 41.6975 0.855 41.7675 0.925 ;
    END
  END rd_sel[12]
  PIN rd_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 45.1625 0.82 45.2325 0.96 ;
      LAYER metal1 ;
        RECT 45.9475 1.2725 46.0825 1.3375 ;
        RECT 45.5875 0.2825 45.6525 0.4175 ;
        RECT 45.165 0.825 45.23 0.96 ;
      LAYER metal2 ;
        RECT 45.9475 1.27 46.0825 1.34 ;
        RECT 45.1625 1.455 46.04 1.525 ;
        RECT 45.97 1.2675 46.04 1.525 ;
        RECT 45.1625 0.4025 45.655 0.4725 ;
        RECT 45.585 0.2825 45.655 0.4725 ;
        RECT 45.1625 0.4025 45.2325 1.525 ;
      LAYER via1 ;
        RECT 45.165 0.86 45.23 0.925 ;
        RECT 45.5875 0.3175 45.6525 0.3825 ;
        RECT 45.9825 1.2725 46.0475 1.3375 ;
      LAYER via2 ;
        RECT 45.1625 0.855 45.2325 0.925 ;
    END
  END rd_sel[13]
  PIN rd_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 48.6275 0.82 48.6975 0.96 ;
      LAYER metal1 ;
        RECT 49.4125 1.2725 49.5475 1.3375 ;
        RECT 49.0525 0.2825 49.1175 0.4175 ;
        RECT 48.63 0.825 48.695 0.96 ;
      LAYER metal2 ;
        RECT 49.4125 1.27 49.5475 1.34 ;
        RECT 48.6275 1.455 49.505 1.525 ;
        RECT 49.435 1.2675 49.505 1.525 ;
        RECT 48.6275 0.4025 49.12 0.4725 ;
        RECT 49.05 0.2825 49.12 0.4725 ;
        RECT 48.6275 0.4025 48.6975 1.525 ;
      LAYER via1 ;
        RECT 48.63 0.86 48.695 0.925 ;
        RECT 49.0525 0.3175 49.1175 0.3825 ;
        RECT 49.4475 1.2725 49.5125 1.3375 ;
      LAYER via2 ;
        RECT 48.6275 0.855 48.6975 0.925 ;
    END
  END rd_sel[14]
  PIN rd_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 52.0925 0.82 52.1625 0.96 ;
      LAYER metal1 ;
        RECT 52.8775 1.2725 53.0125 1.3375 ;
        RECT 52.5175 0.2825 52.5825 0.4175 ;
        RECT 52.095 0.825 52.16 0.96 ;
      LAYER metal2 ;
        RECT 52.8775 1.27 53.0125 1.34 ;
        RECT 52.0925 1.455 52.97 1.525 ;
        RECT 52.9 1.2675 52.97 1.525 ;
        RECT 52.0925 0.4025 52.585 0.4725 ;
        RECT 52.515 0.2825 52.585 0.4725 ;
        RECT 52.0925 0.4025 52.1625 1.525 ;
      LAYER via1 ;
        RECT 52.095 0.86 52.16 0.925 ;
        RECT 52.5175 0.3175 52.5825 0.3825 ;
        RECT 52.9125 1.2725 52.9775 1.3375 ;
      LAYER via2 ;
        RECT 52.0925 0.855 52.1625 0.925 ;
    END
  END rd_sel[15]
  PIN rd_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 55.5575 0.82 55.6275 0.96 ;
      LAYER metal1 ;
        RECT 56.3425 1.2725 56.4775 1.3375 ;
        RECT 55.9825 0.2825 56.0475 0.4175 ;
        RECT 55.56 0.825 55.625 0.96 ;
      LAYER metal2 ;
        RECT 56.3425 1.27 56.4775 1.34 ;
        RECT 55.5575 1.455 56.435 1.525 ;
        RECT 56.365 1.2675 56.435 1.525 ;
        RECT 55.5575 0.4025 56.05 0.4725 ;
        RECT 55.98 0.2825 56.05 0.4725 ;
        RECT 55.5575 0.4025 55.6275 1.525 ;
      LAYER via1 ;
        RECT 55.56 0.86 55.625 0.925 ;
        RECT 55.9825 0.3175 56.0475 0.3825 ;
        RECT 56.3775 1.2725 56.4425 1.3375 ;
      LAYER via2 ;
        RECT 55.5575 0.855 55.6275 0.925 ;
    END
  END rd_sel[16]
  PIN rd_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 59.0225 0.82 59.0925 0.96 ;
      LAYER metal1 ;
        RECT 59.8075 1.2725 59.9425 1.3375 ;
        RECT 59.4475 0.2825 59.5125 0.4175 ;
        RECT 59.025 0.825 59.09 0.96 ;
      LAYER metal2 ;
        RECT 59.8075 1.27 59.9425 1.34 ;
        RECT 59.0225 1.455 59.9 1.525 ;
        RECT 59.83 1.2675 59.9 1.525 ;
        RECT 59.0225 0.4025 59.515 0.4725 ;
        RECT 59.445 0.2825 59.515 0.4725 ;
        RECT 59.0225 0.4025 59.0925 1.525 ;
      LAYER via1 ;
        RECT 59.025 0.86 59.09 0.925 ;
        RECT 59.4475 0.3175 59.5125 0.3825 ;
        RECT 59.8425 1.2725 59.9075 1.3375 ;
      LAYER via2 ;
        RECT 59.0225 0.855 59.0925 0.925 ;
    END
  END rd_sel[17]
  PIN rd_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 62.4875 0.82 62.5575 0.96 ;
      LAYER metal1 ;
        RECT 63.2725 1.2725 63.4075 1.3375 ;
        RECT 62.9125 0.2825 62.9775 0.4175 ;
        RECT 62.49 0.825 62.555 0.96 ;
      LAYER metal2 ;
        RECT 63.2725 1.27 63.4075 1.34 ;
        RECT 62.4875 1.455 63.365 1.525 ;
        RECT 63.295 1.2675 63.365 1.525 ;
        RECT 62.4875 0.4025 62.98 0.4725 ;
        RECT 62.91 0.2825 62.98 0.4725 ;
        RECT 62.4875 0.4025 62.5575 1.525 ;
      LAYER via1 ;
        RECT 62.49 0.86 62.555 0.925 ;
        RECT 62.9125 0.3175 62.9775 0.3825 ;
        RECT 63.3075 1.2725 63.3725 1.3375 ;
      LAYER via2 ;
        RECT 62.4875 0.855 62.5575 0.925 ;
    END
  END rd_sel[18]
  PIN rd_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 65.9525 0.82 66.0225 0.96 ;
      LAYER metal1 ;
        RECT 66.7375 1.2725 66.8725 1.3375 ;
        RECT 66.3775 0.2825 66.4425 0.4175 ;
        RECT 65.955 0.825 66.02 0.96 ;
      LAYER metal2 ;
        RECT 66.7375 1.27 66.8725 1.34 ;
        RECT 65.9525 1.455 66.83 1.525 ;
        RECT 66.76 1.2675 66.83 1.525 ;
        RECT 65.9525 0.4025 66.445 0.4725 ;
        RECT 66.375 0.2825 66.445 0.4725 ;
        RECT 65.9525 0.4025 66.0225 1.525 ;
      LAYER via1 ;
        RECT 65.955 0.86 66.02 0.925 ;
        RECT 66.3775 0.3175 66.4425 0.3825 ;
        RECT 66.7725 1.2725 66.8375 1.3375 ;
      LAYER via2 ;
        RECT 65.9525 0.855 66.0225 0.925 ;
    END
  END rd_sel[19]
  PIN rd_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 3.5825 0.82 3.6525 0.96 ;
      LAYER metal1 ;
        RECT 4.3675 1.2725 4.5025 1.3375 ;
        RECT 4.0075 0.2825 4.0725 0.4175 ;
        RECT 3.585 0.825 3.65 0.96 ;
      LAYER metal2 ;
        RECT 4.3675 1.27 4.5025 1.34 ;
        RECT 3.5825 1.455 4.46 1.525 ;
        RECT 4.39 1.2675 4.46 1.525 ;
        RECT 3.5825 0.4025 4.075 0.4725 ;
        RECT 4.005 0.2825 4.075 0.4725 ;
        RECT 3.5825 0.4025 3.6525 1.525 ;
      LAYER via1 ;
        RECT 3.585 0.86 3.65 0.925 ;
        RECT 4.0075 0.3175 4.0725 0.3825 ;
        RECT 4.4025 1.2725 4.4675 1.3375 ;
      LAYER via2 ;
        RECT 3.5825 0.855 3.6525 0.925 ;
    END
  END rd_sel[1]
  PIN rd_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 69.4175 0.82 69.4875 0.96 ;
      LAYER metal1 ;
        RECT 70.2025 1.2725 70.3375 1.3375 ;
        RECT 69.8425 0.2825 69.9075 0.4175 ;
        RECT 69.42 0.825 69.485 0.96 ;
      LAYER metal2 ;
        RECT 70.2025 1.27 70.3375 1.34 ;
        RECT 69.4175 1.455 70.295 1.525 ;
        RECT 70.225 1.2675 70.295 1.525 ;
        RECT 69.4175 0.4025 69.91 0.4725 ;
        RECT 69.84 0.2825 69.91 0.4725 ;
        RECT 69.4175 0.4025 69.4875 1.525 ;
      LAYER via1 ;
        RECT 69.42 0.86 69.485 0.925 ;
        RECT 69.8425 0.3175 69.9075 0.3825 ;
        RECT 70.2375 1.2725 70.3025 1.3375 ;
      LAYER via2 ;
        RECT 69.4175 0.855 69.4875 0.925 ;
    END
  END rd_sel[20]
  PIN rd_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 72.8825 0.82 72.9525 0.96 ;
      LAYER metal1 ;
        RECT 73.6675 1.2725 73.8025 1.3375 ;
        RECT 73.3075 0.2825 73.3725 0.4175 ;
        RECT 72.885 0.825 72.95 0.96 ;
      LAYER metal2 ;
        RECT 73.6675 1.27 73.8025 1.34 ;
        RECT 72.8825 1.455 73.76 1.525 ;
        RECT 73.69 1.2675 73.76 1.525 ;
        RECT 72.8825 0.4025 73.375 0.4725 ;
        RECT 73.305 0.2825 73.375 0.4725 ;
        RECT 72.8825 0.4025 72.9525 1.525 ;
      LAYER via1 ;
        RECT 72.885 0.86 72.95 0.925 ;
        RECT 73.3075 0.3175 73.3725 0.3825 ;
        RECT 73.7025 1.2725 73.7675 1.3375 ;
      LAYER via2 ;
        RECT 72.8825 0.855 72.9525 0.925 ;
    END
  END rd_sel[21]
  PIN rd_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 76.3475 0.82 76.4175 0.96 ;
      LAYER metal1 ;
        RECT 77.1325 1.2725 77.2675 1.3375 ;
        RECT 76.7725 0.2825 76.8375 0.4175 ;
        RECT 76.35 0.825 76.415 0.96 ;
      LAYER metal2 ;
        RECT 77.1325 1.27 77.2675 1.34 ;
        RECT 76.3475 1.455 77.225 1.525 ;
        RECT 77.155 1.2675 77.225 1.525 ;
        RECT 76.3475 0.4025 76.84 0.4725 ;
        RECT 76.77 0.2825 76.84 0.4725 ;
        RECT 76.3475 0.4025 76.4175 1.525 ;
      LAYER via1 ;
        RECT 76.35 0.86 76.415 0.925 ;
        RECT 76.7725 0.3175 76.8375 0.3825 ;
        RECT 77.1675 1.2725 77.2325 1.3375 ;
      LAYER via2 ;
        RECT 76.3475 0.855 76.4175 0.925 ;
    END
  END rd_sel[22]
  PIN rd_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 79.8125 0.82 79.8825 0.96 ;
      LAYER metal1 ;
        RECT 80.5975 1.2725 80.7325 1.3375 ;
        RECT 80.2375 0.2825 80.3025 0.4175 ;
        RECT 79.815 0.825 79.88 0.96 ;
      LAYER metal2 ;
        RECT 80.5975 1.27 80.7325 1.34 ;
        RECT 79.8125 1.455 80.69 1.525 ;
        RECT 80.62 1.2675 80.69 1.525 ;
        RECT 79.8125 0.4025 80.305 0.4725 ;
        RECT 80.235 0.2825 80.305 0.4725 ;
        RECT 79.8125 0.4025 79.8825 1.525 ;
      LAYER via1 ;
        RECT 79.815 0.86 79.88 0.925 ;
        RECT 80.2375 0.3175 80.3025 0.3825 ;
        RECT 80.6325 1.2725 80.6975 1.3375 ;
      LAYER via2 ;
        RECT 79.8125 0.855 79.8825 0.925 ;
    END
  END rd_sel[23]
  PIN rd_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 83.2775 0.82 83.3475 0.96 ;
      LAYER metal1 ;
        RECT 84.0625 1.2725 84.1975 1.3375 ;
        RECT 83.7025 0.2825 83.7675 0.4175 ;
        RECT 83.28 0.825 83.345 0.96 ;
      LAYER metal2 ;
        RECT 84.0625 1.27 84.1975 1.34 ;
        RECT 83.2775 1.455 84.155 1.525 ;
        RECT 84.085 1.2675 84.155 1.525 ;
        RECT 83.2775 0.4025 83.77 0.4725 ;
        RECT 83.7 0.2825 83.77 0.4725 ;
        RECT 83.2775 0.4025 83.3475 1.525 ;
      LAYER via1 ;
        RECT 83.28 0.86 83.345 0.925 ;
        RECT 83.7025 0.3175 83.7675 0.3825 ;
        RECT 84.0975 1.2725 84.1625 1.3375 ;
      LAYER via2 ;
        RECT 83.2775 0.855 83.3475 0.925 ;
    END
  END rd_sel[24]
  PIN rd_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 86.7425 0.82 86.8125 0.96 ;
      LAYER metal1 ;
        RECT 87.5275 1.2725 87.6625 1.3375 ;
        RECT 87.1675 0.2825 87.2325 0.4175 ;
        RECT 86.745 0.825 86.81 0.96 ;
      LAYER metal2 ;
        RECT 87.5275 1.27 87.6625 1.34 ;
        RECT 86.7425 1.455 87.62 1.525 ;
        RECT 87.55 1.2675 87.62 1.525 ;
        RECT 86.7425 0.4025 87.235 0.4725 ;
        RECT 87.165 0.2825 87.235 0.4725 ;
        RECT 86.7425 0.4025 86.8125 1.525 ;
      LAYER via1 ;
        RECT 86.745 0.86 86.81 0.925 ;
        RECT 87.1675 0.3175 87.2325 0.3825 ;
        RECT 87.5625 1.2725 87.6275 1.3375 ;
      LAYER via2 ;
        RECT 86.7425 0.855 86.8125 0.925 ;
    END
  END rd_sel[25]
  PIN rd_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 90.2075 0.82 90.2775 0.96 ;
      LAYER metal1 ;
        RECT 90.9925 1.2725 91.1275 1.3375 ;
        RECT 90.6325 0.2825 90.6975 0.4175 ;
        RECT 90.21 0.825 90.275 0.96 ;
      LAYER metal2 ;
        RECT 90.9925 1.27 91.1275 1.34 ;
        RECT 90.2075 1.455 91.085 1.525 ;
        RECT 91.015 1.2675 91.085 1.525 ;
        RECT 90.2075 0.4025 90.7 0.4725 ;
        RECT 90.63 0.2825 90.7 0.4725 ;
        RECT 90.2075 0.4025 90.2775 1.525 ;
      LAYER via1 ;
        RECT 90.21 0.86 90.275 0.925 ;
        RECT 90.6325 0.3175 90.6975 0.3825 ;
        RECT 91.0275 1.2725 91.0925 1.3375 ;
      LAYER via2 ;
        RECT 90.2075 0.855 90.2775 0.925 ;
    END
  END rd_sel[26]
  PIN rd_sel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 93.6725 0.82 93.7425 0.96 ;
      LAYER metal1 ;
        RECT 94.4575 1.2725 94.5925 1.3375 ;
        RECT 94.0975 0.2825 94.1625 0.4175 ;
        RECT 93.675 0.825 93.74 0.96 ;
      LAYER metal2 ;
        RECT 94.4575 1.27 94.5925 1.34 ;
        RECT 93.6725 1.455 94.55 1.525 ;
        RECT 94.48 1.2675 94.55 1.525 ;
        RECT 93.6725 0.4025 94.165 0.4725 ;
        RECT 94.095 0.2825 94.165 0.4725 ;
        RECT 93.6725 0.4025 93.7425 1.525 ;
      LAYER via1 ;
        RECT 93.675 0.86 93.74 0.925 ;
        RECT 94.0975 0.3175 94.1625 0.3825 ;
        RECT 94.4925 1.2725 94.5575 1.3375 ;
      LAYER via2 ;
        RECT 93.6725 0.855 93.7425 0.925 ;
    END
  END rd_sel[27]
  PIN rd_sel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 97.1375 0.82 97.2075 0.96 ;
      LAYER metal1 ;
        RECT 97.9225 1.2725 98.0575 1.3375 ;
        RECT 97.5625 0.2825 97.6275 0.4175 ;
        RECT 97.14 0.825 97.205 0.96 ;
      LAYER metal2 ;
        RECT 97.9225 1.27 98.0575 1.34 ;
        RECT 97.1375 1.455 98.015 1.525 ;
        RECT 97.945 1.2675 98.015 1.525 ;
        RECT 97.1375 0.4025 97.63 0.4725 ;
        RECT 97.56 0.2825 97.63 0.4725 ;
        RECT 97.1375 0.4025 97.2075 1.525 ;
      LAYER via1 ;
        RECT 97.14 0.86 97.205 0.925 ;
        RECT 97.5625 0.3175 97.6275 0.3825 ;
        RECT 97.9575 1.2725 98.0225 1.3375 ;
      LAYER via2 ;
        RECT 97.1375 0.855 97.2075 0.925 ;
    END
  END rd_sel[28]
  PIN rd_sel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 100.6025 0.82 100.6725 0.96 ;
      LAYER metal1 ;
        RECT 101.3875 1.2725 101.5225 1.3375 ;
        RECT 101.0275 0.2825 101.0925 0.4175 ;
        RECT 100.605 0.825 100.67 0.96 ;
      LAYER metal2 ;
        RECT 101.3875 1.27 101.5225 1.34 ;
        RECT 100.6025 1.455 101.48 1.525 ;
        RECT 101.41 1.2675 101.48 1.525 ;
        RECT 100.6025 0.4025 101.095 0.4725 ;
        RECT 101.025 0.2825 101.095 0.4725 ;
        RECT 100.6025 0.4025 100.6725 1.525 ;
      LAYER via1 ;
        RECT 100.605 0.86 100.67 0.925 ;
        RECT 101.0275 0.3175 101.0925 0.3825 ;
        RECT 101.4225 1.2725 101.4875 1.3375 ;
      LAYER via2 ;
        RECT 100.6025 0.855 100.6725 0.925 ;
    END
  END rd_sel[29]
  PIN rd_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 7.0475 0.82 7.1175 0.96 ;
      LAYER metal1 ;
        RECT 7.8325 1.2725 7.9675 1.3375 ;
        RECT 7.4725 0.2825 7.5375 0.4175 ;
        RECT 7.05 0.825 7.115 0.96 ;
      LAYER metal2 ;
        RECT 7.8325 1.27 7.9675 1.34 ;
        RECT 7.0475 1.455 7.925 1.525 ;
        RECT 7.855 1.2675 7.925 1.525 ;
        RECT 7.0475 0.4025 7.54 0.4725 ;
        RECT 7.47 0.2825 7.54 0.4725 ;
        RECT 7.0475 0.4025 7.1175 1.525 ;
      LAYER via1 ;
        RECT 7.05 0.86 7.115 0.925 ;
        RECT 7.4725 0.3175 7.5375 0.3825 ;
        RECT 7.8675 1.2725 7.9325 1.3375 ;
      LAYER via2 ;
        RECT 7.0475 0.855 7.1175 0.925 ;
    END
  END rd_sel[2]
  PIN rd_sel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 104.0675 0.82 104.1375 0.96 ;
      LAYER metal1 ;
        RECT 104.8525 1.2725 104.9875 1.3375 ;
        RECT 104.4925 0.2825 104.5575 0.4175 ;
        RECT 104.07 0.825 104.135 0.96 ;
      LAYER metal2 ;
        RECT 104.8525 1.27 104.9875 1.34 ;
        RECT 104.0675 1.455 104.945 1.525 ;
        RECT 104.875 1.2675 104.945 1.525 ;
        RECT 104.0675 0.4025 104.56 0.4725 ;
        RECT 104.49 0.2825 104.56 0.4725 ;
        RECT 104.0675 0.4025 104.1375 1.525 ;
      LAYER via1 ;
        RECT 104.07 0.86 104.135 0.925 ;
        RECT 104.4925 0.3175 104.5575 0.3825 ;
        RECT 104.8875 1.2725 104.9525 1.3375 ;
      LAYER via2 ;
        RECT 104.0675 0.855 104.1375 0.925 ;
    END
  END rd_sel[30]
  PIN rd_sel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 107.5325 0.82 107.6025 0.96 ;
      LAYER metal1 ;
        RECT 108.3175 1.2725 108.4525 1.3375 ;
        RECT 107.9575 0.2825 108.0225 0.4175 ;
        RECT 107.535 0.825 107.6 0.96 ;
      LAYER metal2 ;
        RECT 108.3175 1.27 108.4525 1.34 ;
        RECT 107.5325 1.455 108.41 1.525 ;
        RECT 108.34 1.2675 108.41 1.525 ;
        RECT 107.5325 0.4025 108.025 0.4725 ;
        RECT 107.955 0.2825 108.025 0.4725 ;
        RECT 107.5325 0.4025 107.6025 1.525 ;
      LAYER via1 ;
        RECT 107.535 0.86 107.6 0.925 ;
        RECT 107.9575 0.3175 108.0225 0.3825 ;
        RECT 108.3525 1.2725 108.4175 1.3375 ;
      LAYER via2 ;
        RECT 107.5325 0.855 107.6025 0.925 ;
    END
  END rd_sel[31]
  PIN rd_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 10.5125 0.82 10.5825 0.96 ;
      LAYER metal1 ;
        RECT 11.2975 1.2725 11.4325 1.3375 ;
        RECT 10.9375 0.2825 11.0025 0.4175 ;
        RECT 10.515 0.825 10.58 0.96 ;
      LAYER metal2 ;
        RECT 11.2975 1.27 11.4325 1.34 ;
        RECT 10.5125 1.455 11.39 1.525 ;
        RECT 11.32 1.2675 11.39 1.525 ;
        RECT 10.5125 0.4025 11.005 0.4725 ;
        RECT 10.935 0.2825 11.005 0.4725 ;
        RECT 10.5125 0.4025 10.5825 1.525 ;
      LAYER via1 ;
        RECT 10.515 0.86 10.58 0.925 ;
        RECT 10.9375 0.3175 11.0025 0.3825 ;
        RECT 11.3325 1.2725 11.3975 1.3375 ;
      LAYER via2 ;
        RECT 10.5125 0.855 10.5825 0.925 ;
    END
  END rd_sel[3]
  PIN rd_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 13.9775 0.82 14.0475 0.96 ;
      LAYER metal1 ;
        RECT 14.7625 1.2725 14.8975 1.3375 ;
        RECT 14.4025 0.2825 14.4675 0.4175 ;
        RECT 13.98 0.825 14.045 0.96 ;
      LAYER metal2 ;
        RECT 14.7625 1.27 14.8975 1.34 ;
        RECT 13.9775 1.455 14.855 1.525 ;
        RECT 14.785 1.2675 14.855 1.525 ;
        RECT 13.9775 0.4025 14.47 0.4725 ;
        RECT 14.4 0.2825 14.47 0.4725 ;
        RECT 13.9775 0.4025 14.0475 1.525 ;
      LAYER via1 ;
        RECT 13.98 0.86 14.045 0.925 ;
        RECT 14.4025 0.3175 14.4675 0.3825 ;
        RECT 14.7975 1.2725 14.8625 1.3375 ;
      LAYER via2 ;
        RECT 13.9775 0.855 14.0475 0.925 ;
    END
  END rd_sel[4]
  PIN rd_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 17.4425 0.82 17.5125 0.96 ;
      LAYER metal1 ;
        RECT 18.2275 1.2725 18.3625 1.3375 ;
        RECT 17.8675 0.2825 17.9325 0.4175 ;
        RECT 17.445 0.825 17.51 0.96 ;
      LAYER metal2 ;
        RECT 18.2275 1.27 18.3625 1.34 ;
        RECT 17.4425 1.455 18.32 1.525 ;
        RECT 18.25 1.2675 18.32 1.525 ;
        RECT 17.4425 0.4025 17.935 0.4725 ;
        RECT 17.865 0.2825 17.935 0.4725 ;
        RECT 17.4425 0.4025 17.5125 1.525 ;
      LAYER via1 ;
        RECT 17.445 0.86 17.51 0.925 ;
        RECT 17.8675 0.3175 17.9325 0.3825 ;
        RECT 18.2625 1.2725 18.3275 1.3375 ;
      LAYER via2 ;
        RECT 17.4425 0.855 17.5125 0.925 ;
    END
  END rd_sel[5]
  PIN rd_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 20.9075 0.82 20.9775 0.96 ;
      LAYER metal1 ;
        RECT 21.6925 1.2725 21.8275 1.3375 ;
        RECT 21.3325 0.2825 21.3975 0.4175 ;
        RECT 20.91 0.825 20.975 0.96 ;
      LAYER metal2 ;
        RECT 21.6925 1.27 21.8275 1.34 ;
        RECT 20.9075 1.455 21.785 1.525 ;
        RECT 21.715 1.2675 21.785 1.525 ;
        RECT 20.9075 0.4025 21.4 0.4725 ;
        RECT 21.33 0.2825 21.4 0.4725 ;
        RECT 20.9075 0.4025 20.9775 1.525 ;
      LAYER via1 ;
        RECT 20.91 0.86 20.975 0.925 ;
        RECT 21.3325 0.3175 21.3975 0.3825 ;
        RECT 21.7275 1.2725 21.7925 1.3375 ;
      LAYER via2 ;
        RECT 20.9075 0.855 20.9775 0.925 ;
    END
  END rd_sel[6]
  PIN rd_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 24.3725 0.82 24.4425 0.96 ;
      LAYER metal1 ;
        RECT 25.1575 1.2725 25.2925 1.3375 ;
        RECT 24.7975 0.2825 24.8625 0.4175 ;
        RECT 24.375 0.825 24.44 0.96 ;
      LAYER metal2 ;
        RECT 25.1575 1.27 25.2925 1.34 ;
        RECT 24.3725 1.455 25.25 1.525 ;
        RECT 25.18 1.2675 25.25 1.525 ;
        RECT 24.3725 0.4025 24.865 0.4725 ;
        RECT 24.795 0.2825 24.865 0.4725 ;
        RECT 24.3725 0.4025 24.4425 1.525 ;
      LAYER via1 ;
        RECT 24.375 0.86 24.44 0.925 ;
        RECT 24.7975 0.3175 24.8625 0.3825 ;
        RECT 25.1925 1.2725 25.2575 1.3375 ;
      LAYER via2 ;
        RECT 24.3725 0.855 24.4425 0.925 ;
    END
  END rd_sel[7]
  PIN rd_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 27.8375 0.82 27.9075 0.96 ;
      LAYER metal1 ;
        RECT 28.6225 1.2725 28.7575 1.3375 ;
        RECT 28.2625 0.2825 28.3275 0.4175 ;
        RECT 27.84 0.825 27.905 0.96 ;
      LAYER metal2 ;
        RECT 28.6225 1.27 28.7575 1.34 ;
        RECT 27.8375 1.455 28.715 1.525 ;
        RECT 28.645 1.2675 28.715 1.525 ;
        RECT 27.8375 0.4025 28.33 0.4725 ;
        RECT 28.26 0.2825 28.33 0.4725 ;
        RECT 27.8375 0.4025 27.9075 1.525 ;
      LAYER via1 ;
        RECT 27.84 0.86 27.905 0.925 ;
        RECT 28.2625 0.3175 28.3275 0.3825 ;
        RECT 28.6575 1.2725 28.7225 1.3375 ;
      LAYER via2 ;
        RECT 27.8375 0.855 27.9075 0.925 ;
    END
  END rd_sel[8]
  PIN rd_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 31.3025 0.82 31.3725 0.96 ;
      LAYER metal1 ;
        RECT 32.0875 1.2725 32.2225 1.3375 ;
        RECT 31.7275 0.2825 31.7925 0.4175 ;
        RECT 31.305 0.825 31.37 0.96 ;
      LAYER metal2 ;
        RECT 32.0875 1.27 32.2225 1.34 ;
        RECT 31.3025 1.455 32.18 1.525 ;
        RECT 32.11 1.2675 32.18 1.525 ;
        RECT 31.3025 0.4025 31.795 0.4725 ;
        RECT 31.725 0.2825 31.795 0.4725 ;
        RECT 31.3025 0.4025 31.3725 1.525 ;
      LAYER via1 ;
        RECT 31.305 0.86 31.37 0.925 ;
        RECT 31.7275 0.3175 31.7925 0.3825 ;
        RECT 32.1225 1.2725 32.1875 1.3375 ;
      LAYER via2 ;
        RECT 31.3025 0.855 31.3725 0.925 ;
    END
  END rd_sel[9]
  PIN rd_wdata
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 3.89 1.375 107.91 1.445 ;
        RECT 107.84 0.845 107.91 1.445 ;
        RECT 104.375 0.845 104.445 1.445 ;
        RECT 100.91 0.845 100.98 1.445 ;
        RECT 97.445 0.845 97.515 1.445 ;
        RECT 93.98 0.845 94.05 1.445 ;
        RECT 90.515 0.845 90.585 1.445 ;
        RECT 87.05 0.845 87.12 1.445 ;
        RECT 83.585 0.845 83.655 1.445 ;
        RECT 80.12 0.845 80.19 1.445 ;
        RECT 76.655 0.845 76.725 1.445 ;
        RECT 73.19 0.845 73.26 1.445 ;
        RECT 69.725 0.845 69.795 1.445 ;
        RECT 66.26 0.845 66.33 1.445 ;
        RECT 62.795 0.845 62.865 1.445 ;
        RECT 59.33 0.845 59.4 1.445 ;
        RECT 55.865 0.845 55.935 1.445 ;
        RECT 52.4 0.845 52.47 1.445 ;
        RECT 48.935 0.845 49.005 1.445 ;
        RECT 45.47 0.845 45.54 1.445 ;
        RECT 42.005 0.845 42.075 1.445 ;
        RECT 38.54 0.845 38.61 1.445 ;
        RECT 35.075 0.845 35.145 1.445 ;
        RECT 31.61 0.845 31.68 1.445 ;
        RECT 28.145 0.845 28.215 1.445 ;
        RECT 24.68 0.845 24.75 1.59 ;
        RECT 21.215 0.845 21.285 1.445 ;
        RECT 17.75 0.845 17.82 1.445 ;
        RECT 14.285 0.845 14.355 1.445 ;
        RECT 10.82 0.845 10.89 1.445 ;
        RECT 7.355 0.845 7.425 1.445 ;
        RECT 3.89 0.845 3.96 1.445 ;
      LAYER metal1 ;
        RECT 107.86 0.4875 107.925 1.14 ;
        RECT 107.8425 0.8475 107.925 0.9825 ;
        RECT 104.395 0.4875 104.46 1.14 ;
        RECT 104.3775 0.8475 104.46 0.9825 ;
        RECT 100.93 0.4875 100.995 1.14 ;
        RECT 100.9125 0.8475 100.995 0.9825 ;
        RECT 97.465 0.4875 97.53 1.14 ;
        RECT 97.4475 0.8475 97.53 0.9825 ;
        RECT 94 0.4875 94.065 1.14 ;
        RECT 93.9825 0.8475 94.065 0.9825 ;
        RECT 90.535 0.4875 90.6 1.14 ;
        RECT 90.5175 0.8475 90.6 0.9825 ;
        RECT 87.07 0.4875 87.135 1.14 ;
        RECT 87.0525 0.8475 87.135 0.9825 ;
        RECT 83.605 0.4875 83.67 1.14 ;
        RECT 83.5875 0.8475 83.67 0.9825 ;
        RECT 80.14 0.4875 80.205 1.14 ;
        RECT 80.1225 0.8475 80.205 0.9825 ;
        RECT 76.675 0.4875 76.74 1.14 ;
        RECT 76.6575 0.8475 76.74 0.9825 ;
        RECT 73.21 0.4875 73.275 1.14 ;
        RECT 73.1925 0.8475 73.275 0.9825 ;
        RECT 69.745 0.4875 69.81 1.14 ;
        RECT 69.7275 0.8475 69.81 0.9825 ;
        RECT 66.28 0.4875 66.345 1.14 ;
        RECT 66.2625 0.8475 66.345 0.9825 ;
        RECT 62.815 0.4875 62.88 1.14 ;
        RECT 62.7975 0.8475 62.88 0.9825 ;
        RECT 59.35 0.4875 59.415 1.14 ;
        RECT 59.3325 0.8475 59.415 0.9825 ;
        RECT 55.885 0.4875 55.95 1.14 ;
        RECT 55.8675 0.8475 55.95 0.9825 ;
        RECT 52.42 0.4875 52.485 1.14 ;
        RECT 52.4025 0.8475 52.485 0.9825 ;
        RECT 48.955 0.4875 49.02 1.14 ;
        RECT 48.9375 0.8475 49.02 0.9825 ;
        RECT 45.49 0.4875 45.555 1.14 ;
        RECT 45.4725 0.8475 45.555 0.9825 ;
        RECT 42.025 0.4875 42.09 1.14 ;
        RECT 42.0075 0.8475 42.09 0.9825 ;
        RECT 38.56 0.4875 38.625 1.14 ;
        RECT 38.5425 0.8475 38.625 0.9825 ;
        RECT 35.095 0.4875 35.16 1.14 ;
        RECT 35.0775 0.8475 35.16 0.9825 ;
        RECT 31.63 0.4875 31.695 1.14 ;
        RECT 31.6125 0.8475 31.695 0.9825 ;
        RECT 28.165 0.4875 28.23 1.14 ;
        RECT 28.1475 0.8475 28.23 0.9825 ;
        RECT 24.7 0.4875 24.765 1.14 ;
        RECT 24.6825 0.8475 24.765 0.9825 ;
        RECT 21.235 0.4875 21.3 1.14 ;
        RECT 21.2175 0.8475 21.3 0.9825 ;
        RECT 17.77 0.4875 17.835 1.14 ;
        RECT 17.7525 0.8475 17.835 0.9825 ;
        RECT 14.305 0.4875 14.37 1.14 ;
        RECT 14.2875 0.8475 14.37 0.9825 ;
        RECT 10.84 0.4875 10.905 1.14 ;
        RECT 10.8225 0.8475 10.905 0.9825 ;
        RECT 7.375 0.4875 7.44 1.14 ;
        RECT 7.3575 0.8475 7.44 0.9825 ;
        RECT 3.91 0.4875 3.975 1.14 ;
        RECT 3.8925 0.8475 3.975 0.9825 ;
      LAYER metal2 ;
        RECT 107.84 0.845 107.91 0.985 ;
        RECT 104.375 0.845 104.445 0.985 ;
        RECT 100.91 0.845 100.98 0.985 ;
        RECT 97.445 0.845 97.515 0.985 ;
        RECT 93.98 0.845 94.05 0.985 ;
        RECT 90.515 0.845 90.585 0.985 ;
        RECT 87.05 0.845 87.12 0.985 ;
        RECT 83.585 0.845 83.655 0.985 ;
        RECT 80.12 0.845 80.19 0.985 ;
        RECT 76.655 0.845 76.725 0.985 ;
        RECT 73.19 0.845 73.26 0.985 ;
        RECT 69.725 0.845 69.795 0.985 ;
        RECT 66.26 0.845 66.33 0.985 ;
        RECT 62.795 0.845 62.865 0.985 ;
        RECT 59.33 0.845 59.4 0.985 ;
        RECT 55.865 0.845 55.935 0.985 ;
        RECT 52.4 0.845 52.47 0.985 ;
        RECT 48.935 0.845 49.005 0.985 ;
        RECT 45.47 0.845 45.54 0.985 ;
        RECT 42.005 0.845 42.075 0.985 ;
        RECT 38.54 0.845 38.61 0.985 ;
        RECT 35.075 0.845 35.145 0.985 ;
        RECT 31.61 0.845 31.68 0.985 ;
        RECT 28.145 0.845 28.215 0.985 ;
        RECT 24.68 0.845 24.75 0.985 ;
        RECT 21.215 0.845 21.285 0.985 ;
        RECT 17.75 0.845 17.82 0.985 ;
        RECT 14.285 0.845 14.355 0.985 ;
        RECT 10.82 0.845 10.89 0.985 ;
        RECT 7.355 0.845 7.425 0.985 ;
        RECT 3.89 0.845 3.96 0.985 ;
      LAYER via1 ;
        RECT 3.8925 0.8825 3.9575 0.9475 ;
        RECT 7.3575 0.8825 7.4225 0.9475 ;
        RECT 10.8225 0.8825 10.8875 0.9475 ;
        RECT 14.2875 0.8825 14.3525 0.9475 ;
        RECT 17.7525 0.8825 17.8175 0.9475 ;
        RECT 21.2175 0.8825 21.2825 0.9475 ;
        RECT 24.6825 0.8825 24.7475 0.9475 ;
        RECT 28.1475 0.8825 28.2125 0.9475 ;
        RECT 31.6125 0.8825 31.6775 0.9475 ;
        RECT 35.0775 0.8825 35.1425 0.9475 ;
        RECT 38.5425 0.8825 38.6075 0.9475 ;
        RECT 42.0075 0.8825 42.0725 0.9475 ;
        RECT 45.4725 0.8825 45.5375 0.9475 ;
        RECT 48.9375 0.8825 49.0025 0.9475 ;
        RECT 52.4025 0.8825 52.4675 0.9475 ;
        RECT 55.8675 0.8825 55.9325 0.9475 ;
        RECT 59.3325 0.8825 59.3975 0.9475 ;
        RECT 62.7975 0.8825 62.8625 0.9475 ;
        RECT 66.2625 0.8825 66.3275 0.9475 ;
        RECT 69.7275 0.8825 69.7925 0.9475 ;
        RECT 73.1925 0.8825 73.2575 0.9475 ;
        RECT 76.6575 0.8825 76.7225 0.9475 ;
        RECT 80.1225 0.8825 80.1875 0.9475 ;
        RECT 83.5875 0.8825 83.6525 0.9475 ;
        RECT 87.0525 0.8825 87.1175 0.9475 ;
        RECT 90.5175 0.8825 90.5825 0.9475 ;
        RECT 93.9825 0.8825 94.0475 0.9475 ;
        RECT 97.4475 0.8825 97.5125 0.9475 ;
        RECT 100.9125 0.8825 100.9775 0.9475 ;
        RECT 104.3775 0.8825 104.4425 0.9475 ;
        RECT 107.8425 0.8825 107.9075 0.9475 ;
      LAYER via2 ;
        RECT 3.89 0.88 3.96 0.95 ;
        RECT 7.355 0.88 7.425 0.95 ;
        RECT 10.82 0.88 10.89 0.95 ;
        RECT 14.285 0.88 14.355 0.95 ;
        RECT 17.75 0.88 17.82 0.95 ;
        RECT 21.215 0.88 21.285 0.95 ;
        RECT 24.68 0.88 24.75 0.95 ;
        RECT 28.145 0.88 28.215 0.95 ;
        RECT 31.61 0.88 31.68 0.95 ;
        RECT 35.075 0.88 35.145 0.95 ;
        RECT 38.54 0.88 38.61 0.95 ;
        RECT 42.005 0.88 42.075 0.95 ;
        RECT 45.47 0.88 45.54 0.95 ;
        RECT 48.935 0.88 49.005 0.95 ;
        RECT 52.4 0.88 52.47 0.95 ;
        RECT 55.865 0.88 55.935 0.95 ;
        RECT 59.33 0.88 59.4 0.95 ;
        RECT 62.795 0.88 62.865 0.95 ;
        RECT 66.26 0.88 66.33 0.95 ;
        RECT 69.725 0.88 69.795 0.95 ;
        RECT 73.19 0.88 73.26 0.95 ;
        RECT 76.655 0.88 76.725 0.95 ;
        RECT 80.12 0.88 80.19 0.95 ;
        RECT 83.585 0.88 83.655 0.95 ;
        RECT 87.05 0.88 87.12 0.95 ;
        RECT 90.515 0.88 90.585 0.95 ;
        RECT 93.98 0.88 94.05 0.95 ;
        RECT 97.445 0.88 97.515 0.95 ;
        RECT 100.91 0.88 100.98 0.95 ;
        RECT 104.375 0.88 104.445 0.95 ;
        RECT 107.84 0.88 107.91 0.95 ;
    END
  END rd_wdata
  PIN rs1_rdata
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 112.045 1.03 112.11 1.165 ;
        RECT 111.71 0.265 111.775 1.355 ;
      LAYER metal2 ;
        RECT 112.04 1.03 112.1125 1.165 ;
        RECT 112.04 0.89 112.11 1.165 ;
        RECT 111.7075 0.89 112.11 0.96 ;
        RECT 111.7075 0.89 111.7775 1.355 ;
      LAYER via1 ;
        RECT 111.71 1.255 111.775 1.32 ;
        RECT 112.045 1.065 112.11 1.13 ;
    END
  END rs1_rdata
  PIN rs1_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.28 0.455 3.345 0.59 ;
        RECT 2.0875 0.265 2.1525 0.4 ;
      LAYER metal2 ;
        RECT 3.2775 0.125 3.3475 0.59 ;
        RECT 2.0825 0.125 3.3475 0.195 ;
        RECT 2.0825 0.265 2.155 0.4 ;
        RECT 2.0825 0.125 2.1525 0.4 ;
      LAYER via1 ;
        RECT 2.0875 0.3 2.1525 0.365 ;
        RECT 3.28 0.49 3.345 0.555 ;
    END
  END rs1_sel[0]
  PIN rs1_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 37.93 0.455 37.995 0.59 ;
        RECT 36.7375 0.265 36.8025 0.4 ;
      LAYER metal2 ;
        RECT 37.9275 0.125 37.9975 0.59 ;
        RECT 36.7325 0.125 37.9975 0.195 ;
        RECT 36.7325 0.265 36.805 0.4 ;
        RECT 36.7325 0.125 36.8025 0.4 ;
      LAYER via1 ;
        RECT 36.7375 0.3 36.8025 0.365 ;
        RECT 37.93 0.49 37.995 0.555 ;
    END
  END rs1_sel[10]
  PIN rs1_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 41.395 0.455 41.46 0.59 ;
        RECT 40.2025 0.265 40.2675 0.4 ;
      LAYER metal2 ;
        RECT 41.3925 0.125 41.4625 0.59 ;
        RECT 40.1975 0.125 41.4625 0.195 ;
        RECT 40.1975 0.265 40.27 0.4 ;
        RECT 40.1975 0.125 40.2675 0.4 ;
      LAYER via1 ;
        RECT 40.2025 0.3 40.2675 0.365 ;
        RECT 41.395 0.49 41.46 0.555 ;
    END
  END rs1_sel[11]
  PIN rs1_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 44.86 0.455 44.925 0.59 ;
        RECT 43.6675 0.265 43.7325 0.4 ;
      LAYER metal2 ;
        RECT 44.8575 0.125 44.9275 0.59 ;
        RECT 43.6625 0.125 44.9275 0.195 ;
        RECT 43.6625 0.265 43.735 0.4 ;
        RECT 43.6625 0.125 43.7325 0.4 ;
      LAYER via1 ;
        RECT 43.6675 0.3 43.7325 0.365 ;
        RECT 44.86 0.49 44.925 0.555 ;
    END
  END rs1_sel[12]
  PIN rs1_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 48.325 0.455 48.39 0.59 ;
        RECT 47.1325 0.265 47.1975 0.4 ;
      LAYER metal2 ;
        RECT 48.3225 0.125 48.3925 0.59 ;
        RECT 47.1275 0.125 48.3925 0.195 ;
        RECT 47.1275 0.265 47.2 0.4 ;
        RECT 47.1275 0.125 47.1975 0.4 ;
      LAYER via1 ;
        RECT 47.1325 0.3 47.1975 0.365 ;
        RECT 48.325 0.49 48.39 0.555 ;
    END
  END rs1_sel[13]
  PIN rs1_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 51.79 0.455 51.855 0.59 ;
        RECT 50.5975 0.265 50.6625 0.4 ;
      LAYER metal2 ;
        RECT 51.7875 0.125 51.8575 0.59 ;
        RECT 50.5925 0.125 51.8575 0.195 ;
        RECT 50.5925 0.265 50.665 0.4 ;
        RECT 50.5925 0.125 50.6625 0.4 ;
      LAYER via1 ;
        RECT 50.5975 0.3 50.6625 0.365 ;
        RECT 51.79 0.49 51.855 0.555 ;
    END
  END rs1_sel[14]
  PIN rs1_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 55.255 0.455 55.32 0.59 ;
        RECT 54.0625 0.265 54.1275 0.4 ;
      LAYER metal2 ;
        RECT 55.2525 0.125 55.3225 0.59 ;
        RECT 54.0575 0.125 55.3225 0.195 ;
        RECT 54.0575 0.265 54.13 0.4 ;
        RECT 54.0575 0.125 54.1275 0.4 ;
      LAYER via1 ;
        RECT 54.0625 0.3 54.1275 0.365 ;
        RECT 55.255 0.49 55.32 0.555 ;
    END
  END rs1_sel[15]
  PIN rs1_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 58.72 0.455 58.785 0.59 ;
        RECT 57.5275 0.265 57.5925 0.4 ;
      LAYER metal2 ;
        RECT 58.7175 0.125 58.7875 0.59 ;
        RECT 57.5225 0.125 58.7875 0.195 ;
        RECT 57.5225 0.265 57.595 0.4 ;
        RECT 57.5225 0.125 57.5925 0.4 ;
      LAYER via1 ;
        RECT 57.5275 0.3 57.5925 0.365 ;
        RECT 58.72 0.49 58.785 0.555 ;
    END
  END rs1_sel[16]
  PIN rs1_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 62.185 0.455 62.25 0.59 ;
        RECT 60.9925 0.265 61.0575 0.4 ;
      LAYER metal2 ;
        RECT 62.1825 0.125 62.2525 0.59 ;
        RECT 60.9875 0.125 62.2525 0.195 ;
        RECT 60.9875 0.265 61.06 0.4 ;
        RECT 60.9875 0.125 61.0575 0.4 ;
      LAYER via1 ;
        RECT 60.9925 0.3 61.0575 0.365 ;
        RECT 62.185 0.49 62.25 0.555 ;
    END
  END rs1_sel[17]
  PIN rs1_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 65.65 0.455 65.715 0.59 ;
        RECT 64.4575 0.265 64.5225 0.4 ;
      LAYER metal2 ;
        RECT 65.6475 0.125 65.7175 0.59 ;
        RECT 64.4525 0.125 65.7175 0.195 ;
        RECT 64.4525 0.265 64.525 0.4 ;
        RECT 64.4525 0.125 64.5225 0.4 ;
      LAYER via1 ;
        RECT 64.4575 0.3 64.5225 0.365 ;
        RECT 65.65 0.49 65.715 0.555 ;
    END
  END rs1_sel[18]
  PIN rs1_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 69.115 0.455 69.18 0.59 ;
        RECT 67.9225 0.265 67.9875 0.4 ;
      LAYER metal2 ;
        RECT 69.1125 0.125 69.1825 0.59 ;
        RECT 67.9175 0.125 69.1825 0.195 ;
        RECT 67.9175 0.265 67.99 0.4 ;
        RECT 67.9175 0.125 67.9875 0.4 ;
      LAYER via1 ;
        RECT 67.9225 0.3 67.9875 0.365 ;
        RECT 69.115 0.49 69.18 0.555 ;
    END
  END rs1_sel[19]
  PIN rs1_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.745 0.455 6.81 0.59 ;
        RECT 5.5525 0.265 5.6175 0.4 ;
      LAYER metal2 ;
        RECT 6.7425 0.125 6.8125 0.59 ;
        RECT 5.5475 0.125 6.8125 0.195 ;
        RECT 5.5475 0.265 5.62 0.4 ;
        RECT 5.5475 0.125 5.6175 0.4 ;
      LAYER via1 ;
        RECT 5.5525 0.3 5.6175 0.365 ;
        RECT 6.745 0.49 6.81 0.555 ;
    END
  END rs1_sel[1]
  PIN rs1_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 72.58 0.455 72.645 0.59 ;
        RECT 71.3875 0.265 71.4525 0.4 ;
      LAYER metal2 ;
        RECT 72.5775 0.125 72.6475 0.59 ;
        RECT 71.3825 0.125 72.6475 0.195 ;
        RECT 71.3825 0.265 71.455 0.4 ;
        RECT 71.3825 0.125 71.4525 0.4 ;
      LAYER via1 ;
        RECT 71.3875 0.3 71.4525 0.365 ;
        RECT 72.58 0.49 72.645 0.555 ;
    END
  END rs1_sel[20]
  PIN rs1_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 76.045 0.455 76.11 0.59 ;
        RECT 74.8525 0.265 74.9175 0.4 ;
      LAYER metal2 ;
        RECT 76.0425 0.125 76.1125 0.59 ;
        RECT 74.8475 0.125 76.1125 0.195 ;
        RECT 74.8475 0.265 74.92 0.4 ;
        RECT 74.8475 0.125 74.9175 0.4 ;
      LAYER via1 ;
        RECT 74.8525 0.3 74.9175 0.365 ;
        RECT 76.045 0.49 76.11 0.555 ;
    END
  END rs1_sel[21]
  PIN rs1_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 79.51 0.455 79.575 0.59 ;
        RECT 78.3175 0.265 78.3825 0.4 ;
      LAYER metal2 ;
        RECT 79.5075 0.125 79.5775 0.59 ;
        RECT 78.3125 0.125 79.5775 0.195 ;
        RECT 78.3125 0.265 78.385 0.4 ;
        RECT 78.3125 0.125 78.3825 0.4 ;
      LAYER via1 ;
        RECT 78.3175 0.3 78.3825 0.365 ;
        RECT 79.51 0.49 79.575 0.555 ;
    END
  END rs1_sel[22]
  PIN rs1_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 82.975 0.455 83.04 0.59 ;
        RECT 81.7825 0.265 81.8475 0.4 ;
      LAYER metal2 ;
        RECT 82.9725 0.125 83.0425 0.59 ;
        RECT 81.7775 0.125 83.0425 0.195 ;
        RECT 81.7775 0.265 81.85 0.4 ;
        RECT 81.7775 0.125 81.8475 0.4 ;
      LAYER via1 ;
        RECT 81.7825 0.3 81.8475 0.365 ;
        RECT 82.975 0.49 83.04 0.555 ;
    END
  END rs1_sel[23]
  PIN rs1_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 86.44 0.455 86.505 0.59 ;
        RECT 85.2475 0.265 85.3125 0.4 ;
      LAYER metal2 ;
        RECT 86.4375 0.125 86.5075 0.59 ;
        RECT 85.2425 0.125 86.5075 0.195 ;
        RECT 85.2425 0.265 85.315 0.4 ;
        RECT 85.2425 0.125 85.3125 0.4 ;
      LAYER via1 ;
        RECT 85.2475 0.3 85.3125 0.365 ;
        RECT 86.44 0.49 86.505 0.555 ;
    END
  END rs1_sel[24]
  PIN rs1_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 89.905 0.455 89.97 0.59 ;
        RECT 88.7125 0.265 88.7775 0.4 ;
      LAYER metal2 ;
        RECT 89.9025 0.125 89.9725 0.59 ;
        RECT 88.7075 0.125 89.9725 0.195 ;
        RECT 88.7075 0.265 88.78 0.4 ;
        RECT 88.7075 0.125 88.7775 0.4 ;
      LAYER via1 ;
        RECT 88.7125 0.3 88.7775 0.365 ;
        RECT 89.905 0.49 89.97 0.555 ;
    END
  END rs1_sel[25]
  PIN rs1_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 93.37 0.455 93.435 0.59 ;
        RECT 92.1775 0.265 92.2425 0.4 ;
      LAYER metal2 ;
        RECT 93.3675 0.125 93.4375 0.59 ;
        RECT 92.1725 0.125 93.4375 0.195 ;
        RECT 92.1725 0.265 92.245 0.4 ;
        RECT 92.1725 0.125 92.2425 0.4 ;
      LAYER via1 ;
        RECT 92.1775 0.3 92.2425 0.365 ;
        RECT 93.37 0.49 93.435 0.555 ;
    END
  END rs1_sel[26]
  PIN rs1_sel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 96.835 0.455 96.9 0.59 ;
        RECT 95.6425 0.265 95.7075 0.4 ;
      LAYER metal2 ;
        RECT 96.8325 0.125 96.9025 0.59 ;
        RECT 95.6375 0.125 96.9025 0.195 ;
        RECT 95.6375 0.265 95.71 0.4 ;
        RECT 95.6375 0.125 95.7075 0.4 ;
      LAYER via1 ;
        RECT 95.6425 0.3 95.7075 0.365 ;
        RECT 96.835 0.49 96.9 0.555 ;
    END
  END rs1_sel[27]
  PIN rs1_sel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 100.3 0.455 100.365 0.59 ;
        RECT 99.1075 0.265 99.1725 0.4 ;
      LAYER metal2 ;
        RECT 100.2975 0.125 100.3675 0.59 ;
        RECT 99.1025 0.125 100.3675 0.195 ;
        RECT 99.1025 0.265 99.175 0.4 ;
        RECT 99.1025 0.125 99.1725 0.4 ;
      LAYER via1 ;
        RECT 99.1075 0.3 99.1725 0.365 ;
        RECT 100.3 0.49 100.365 0.555 ;
    END
  END rs1_sel[28]
  PIN rs1_sel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 103.765 0.455 103.83 0.59 ;
        RECT 102.5725 0.265 102.6375 0.4 ;
      LAYER metal2 ;
        RECT 103.7625 0.125 103.8325 0.59 ;
        RECT 102.5675 0.125 103.8325 0.195 ;
        RECT 102.5675 0.265 102.64 0.4 ;
        RECT 102.5675 0.125 102.6375 0.4 ;
      LAYER via1 ;
        RECT 102.5725 0.3 102.6375 0.365 ;
        RECT 103.765 0.49 103.83 0.555 ;
    END
  END rs1_sel[29]
  PIN rs1_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 10.21 0.455 10.275 0.59 ;
        RECT 9.0175 0.265 9.0825 0.4 ;
      LAYER metal2 ;
        RECT 10.2075 0.125 10.2775 0.59 ;
        RECT 9.0125 0.125 10.2775 0.195 ;
        RECT 9.0125 0.265 9.085 0.4 ;
        RECT 9.0125 0.125 9.0825 0.4 ;
      LAYER via1 ;
        RECT 9.0175 0.3 9.0825 0.365 ;
        RECT 10.21 0.49 10.275 0.555 ;
    END
  END rs1_sel[2]
  PIN rs1_sel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 107.23 0.455 107.295 0.59 ;
        RECT 106.0375 0.265 106.1025 0.4 ;
      LAYER metal2 ;
        RECT 107.2275 0.125 107.2975 0.59 ;
        RECT 106.0325 0.125 107.2975 0.195 ;
        RECT 106.0325 0.265 106.105 0.4 ;
        RECT 106.0325 0.125 106.1025 0.4 ;
      LAYER via1 ;
        RECT 106.0375 0.3 106.1025 0.365 ;
        RECT 107.23 0.49 107.295 0.555 ;
    END
  END rs1_sel[30]
  PIN rs1_sel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 110.695 0.455 110.76 0.59 ;
        RECT 109.5025 0.265 109.5675 0.4 ;
      LAYER metal2 ;
        RECT 110.6925 0.125 110.7625 0.59 ;
        RECT 109.4975 0.125 110.7625 0.195 ;
        RECT 109.4975 0.265 109.57 0.4 ;
        RECT 109.4975 0.125 109.5675 0.4 ;
      LAYER via1 ;
        RECT 109.5025 0.3 109.5675 0.365 ;
        RECT 110.695 0.49 110.76 0.555 ;
    END
  END rs1_sel[31]
  PIN rs1_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 13.675 0.455 13.74 0.59 ;
        RECT 12.4825 0.265 12.5475 0.4 ;
      LAYER metal2 ;
        RECT 13.6725 0.125 13.7425 0.59 ;
        RECT 12.4775 0.125 13.7425 0.195 ;
        RECT 12.4775 0.265 12.55 0.4 ;
        RECT 12.4775 0.125 12.5475 0.4 ;
      LAYER via1 ;
        RECT 12.4825 0.3 12.5475 0.365 ;
        RECT 13.675 0.49 13.74 0.555 ;
    END
  END rs1_sel[3]
  PIN rs1_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 17.14 0.455 17.205 0.59 ;
        RECT 15.9475 0.265 16.0125 0.4 ;
      LAYER metal2 ;
        RECT 17.1375 0.125 17.2075 0.59 ;
        RECT 15.9425 0.125 17.2075 0.195 ;
        RECT 15.9425 0.265 16.015 0.4 ;
        RECT 15.9425 0.125 16.0125 0.4 ;
      LAYER via1 ;
        RECT 15.9475 0.3 16.0125 0.365 ;
        RECT 17.14 0.49 17.205 0.555 ;
    END
  END rs1_sel[4]
  PIN rs1_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 20.605 0.455 20.67 0.59 ;
        RECT 19.4125 0.265 19.4775 0.4 ;
      LAYER metal2 ;
        RECT 20.6025 0.125 20.6725 0.59 ;
        RECT 19.4075 0.125 20.6725 0.195 ;
        RECT 19.4075 0.265 19.48 0.4 ;
        RECT 19.4075 0.125 19.4775 0.4 ;
      LAYER via1 ;
        RECT 19.4125 0.3 19.4775 0.365 ;
        RECT 20.605 0.49 20.67 0.555 ;
    END
  END rs1_sel[5]
  PIN rs1_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 24.07 0.455 24.135 0.59 ;
        RECT 22.8775 0.265 22.9425 0.4 ;
      LAYER metal2 ;
        RECT 24.0675 0.125 24.1375 0.59 ;
        RECT 22.8725 0.125 24.1375 0.195 ;
        RECT 22.8725 0.265 22.945 0.4 ;
        RECT 22.8725 0.125 22.9425 0.4 ;
      LAYER via1 ;
        RECT 22.8775 0.3 22.9425 0.365 ;
        RECT 24.07 0.49 24.135 0.555 ;
    END
  END rs1_sel[6]
  PIN rs1_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 27.535 0.455 27.6 0.59 ;
        RECT 26.3425 0.265 26.4075 0.4 ;
      LAYER metal2 ;
        RECT 27.5325 0.125 27.6025 0.59 ;
        RECT 26.3375 0.125 27.6025 0.195 ;
        RECT 26.3375 0.265 26.41 0.4 ;
        RECT 26.3375 0.125 26.4075 0.4 ;
      LAYER via1 ;
        RECT 26.3425 0.3 26.4075 0.365 ;
        RECT 27.535 0.49 27.6 0.555 ;
    END
  END rs1_sel[7]
  PIN rs1_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 31 0.455 31.065 0.59 ;
        RECT 29.8075 0.265 29.8725 0.4 ;
      LAYER metal2 ;
        RECT 30.9975 0.125 31.0675 0.59 ;
        RECT 29.8025 0.125 31.0675 0.195 ;
        RECT 29.8025 0.265 29.875 0.4 ;
        RECT 29.8025 0.125 29.8725 0.4 ;
      LAYER via1 ;
        RECT 29.8075 0.3 29.8725 0.365 ;
        RECT 31 0.49 31.065 0.555 ;
    END
  END rs1_sel[8]
  PIN rs1_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 34.465 0.455 34.53 0.59 ;
        RECT 33.2725 0.265 33.3375 0.4 ;
      LAYER metal2 ;
        RECT 34.4625 0.125 34.5325 0.59 ;
        RECT 33.2675 0.125 34.5325 0.195 ;
        RECT 33.2675 0.265 33.34 0.4 ;
        RECT 33.2675 0.125 33.3375 0.4 ;
      LAYER via1 ;
        RECT 33.2725 0.3 33.3375 0.365 ;
        RECT 34.465 0.49 34.53 0.555 ;
    END
  END rs1_sel[9]
  PIN rs2_rdata
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 115.31 0.265 115.375 1.355 ;
        RECT 114.975 1.03 115.04 1.165 ;
      LAYER metal2 ;
        RECT 115.3075 0.89 115.3775 1.355 ;
        RECT 114.975 0.89 115.3775 0.96 ;
        RECT 114.9725 1.03 115.045 1.165 ;
        RECT 114.975 0.89 115.045 1.165 ;
      LAYER via1 ;
        RECT 114.975 1.065 115.04 1.13 ;
        RECT 115.31 1.255 115.375 1.32 ;
    END
  END rs2_rdata
  PIN rs2_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 2.9175 0.8225 2.9875 0.9625 ;
      LAYER metal1 ;
        RECT 2.9225 0.825 2.9875 0.96 ;
        RECT 2.4675 0.2825 2.5325 0.4175 ;
      LAYER metal2 ;
        RECT 2.9175 0.825 2.99 0.96 ;
        RECT 2.9175 0.315 2.9875 0.9625 ;
        RECT 2.465 0.315 2.9875 0.385 ;
        RECT 2.465 0.2825 2.535 0.4175 ;
      LAYER via1 ;
        RECT 2.4675 0.3175 2.5325 0.3825 ;
        RECT 2.9225 0.86 2.9875 0.925 ;
      LAYER via2 ;
        RECT 2.9175 0.8575 2.9875 0.9275 ;
    END
  END rs2_sel[0]
  PIN rs2_sel[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 37.5675 0.8225 37.6375 0.9625 ;
      LAYER metal1 ;
        RECT 37.5725 0.825 37.6375 0.96 ;
        RECT 37.1175 0.2825 37.1825 0.4175 ;
      LAYER metal2 ;
        RECT 37.5675 0.825 37.64 0.96 ;
        RECT 37.5675 0.315 37.6375 0.9625 ;
        RECT 37.115 0.315 37.6375 0.385 ;
        RECT 37.115 0.2825 37.185 0.4175 ;
      LAYER via1 ;
        RECT 37.1175 0.3175 37.1825 0.3825 ;
        RECT 37.5725 0.86 37.6375 0.925 ;
      LAYER via2 ;
        RECT 37.5675 0.8575 37.6375 0.9275 ;
    END
  END rs2_sel[10]
  PIN rs2_sel[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 41.0325 0.8225 41.1025 0.9625 ;
      LAYER metal1 ;
        RECT 41.0375 0.825 41.1025 0.96 ;
        RECT 40.5825 0.2825 40.6475 0.4175 ;
      LAYER metal2 ;
        RECT 41.0325 0.825 41.105 0.96 ;
        RECT 41.0325 0.315 41.1025 0.9625 ;
        RECT 40.58 0.315 41.1025 0.385 ;
        RECT 40.58 0.2825 40.65 0.4175 ;
      LAYER via1 ;
        RECT 40.5825 0.3175 40.6475 0.3825 ;
        RECT 41.0375 0.86 41.1025 0.925 ;
      LAYER via2 ;
        RECT 41.0325 0.8575 41.1025 0.9275 ;
    END
  END rs2_sel[11]
  PIN rs2_sel[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 44.4975 0.8225 44.5675 0.9625 ;
      LAYER metal1 ;
        RECT 44.5025 0.825 44.5675 0.96 ;
        RECT 44.0475 0.2825 44.1125 0.4175 ;
      LAYER metal2 ;
        RECT 44.4975 0.825 44.57 0.96 ;
        RECT 44.4975 0.315 44.5675 0.9625 ;
        RECT 44.045 0.315 44.5675 0.385 ;
        RECT 44.045 0.2825 44.115 0.4175 ;
      LAYER via1 ;
        RECT 44.0475 0.3175 44.1125 0.3825 ;
        RECT 44.5025 0.86 44.5675 0.925 ;
      LAYER via2 ;
        RECT 44.4975 0.8575 44.5675 0.9275 ;
    END
  END rs2_sel[12]
  PIN rs2_sel[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 47.9625 0.8225 48.0325 0.9625 ;
      LAYER metal1 ;
        RECT 47.9675 0.825 48.0325 0.96 ;
        RECT 47.5125 0.2825 47.5775 0.4175 ;
      LAYER metal2 ;
        RECT 47.9625 0.825 48.035 0.96 ;
        RECT 47.9625 0.315 48.0325 0.9625 ;
        RECT 47.51 0.315 48.0325 0.385 ;
        RECT 47.51 0.2825 47.58 0.4175 ;
      LAYER via1 ;
        RECT 47.5125 0.3175 47.5775 0.3825 ;
        RECT 47.9675 0.86 48.0325 0.925 ;
      LAYER via2 ;
        RECT 47.9625 0.8575 48.0325 0.9275 ;
    END
  END rs2_sel[13]
  PIN rs2_sel[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 51.4275 0.8225 51.4975 0.9625 ;
      LAYER metal1 ;
        RECT 51.4325 0.825 51.4975 0.96 ;
        RECT 50.9775 0.2825 51.0425 0.4175 ;
      LAYER metal2 ;
        RECT 51.4275 0.825 51.5 0.96 ;
        RECT 51.4275 0.315 51.4975 0.9625 ;
        RECT 50.975 0.315 51.4975 0.385 ;
        RECT 50.975 0.2825 51.045 0.4175 ;
      LAYER via1 ;
        RECT 50.9775 0.3175 51.0425 0.3825 ;
        RECT 51.4325 0.86 51.4975 0.925 ;
      LAYER via2 ;
        RECT 51.4275 0.8575 51.4975 0.9275 ;
    END
  END rs2_sel[14]
  PIN rs2_sel[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 54.8925 0.8225 54.9625 0.9625 ;
      LAYER metal1 ;
        RECT 54.8975 0.825 54.9625 0.96 ;
        RECT 54.4425 0.2825 54.5075 0.4175 ;
      LAYER metal2 ;
        RECT 54.8925 0.825 54.965 0.96 ;
        RECT 54.8925 0.315 54.9625 0.9625 ;
        RECT 54.44 0.315 54.9625 0.385 ;
        RECT 54.44 0.2825 54.51 0.4175 ;
      LAYER via1 ;
        RECT 54.4425 0.3175 54.5075 0.3825 ;
        RECT 54.8975 0.86 54.9625 0.925 ;
      LAYER via2 ;
        RECT 54.8925 0.8575 54.9625 0.9275 ;
    END
  END rs2_sel[15]
  PIN rs2_sel[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 58.3575 0.8225 58.4275 0.9625 ;
      LAYER metal1 ;
        RECT 58.3625 0.825 58.4275 0.96 ;
        RECT 57.9075 0.2825 57.9725 0.4175 ;
      LAYER metal2 ;
        RECT 58.3575 0.825 58.43 0.96 ;
        RECT 58.3575 0.315 58.4275 0.9625 ;
        RECT 57.905 0.315 58.4275 0.385 ;
        RECT 57.905 0.2825 57.975 0.4175 ;
      LAYER via1 ;
        RECT 57.9075 0.3175 57.9725 0.3825 ;
        RECT 58.3625 0.86 58.4275 0.925 ;
      LAYER via2 ;
        RECT 58.3575 0.8575 58.4275 0.9275 ;
    END
  END rs2_sel[16]
  PIN rs2_sel[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 61.8225 0.8225 61.8925 0.9625 ;
      LAYER metal1 ;
        RECT 61.8275 0.825 61.8925 0.96 ;
        RECT 61.3725 0.2825 61.4375 0.4175 ;
      LAYER metal2 ;
        RECT 61.8225 0.825 61.895 0.96 ;
        RECT 61.8225 0.315 61.8925 0.9625 ;
        RECT 61.37 0.315 61.8925 0.385 ;
        RECT 61.37 0.2825 61.44 0.4175 ;
      LAYER via1 ;
        RECT 61.3725 0.3175 61.4375 0.3825 ;
        RECT 61.8275 0.86 61.8925 0.925 ;
      LAYER via2 ;
        RECT 61.8225 0.8575 61.8925 0.9275 ;
    END
  END rs2_sel[17]
  PIN rs2_sel[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 65.2875 0.8225 65.3575 0.9625 ;
      LAYER metal1 ;
        RECT 65.2925 0.825 65.3575 0.96 ;
        RECT 64.8375 0.2825 64.9025 0.4175 ;
      LAYER metal2 ;
        RECT 65.2875 0.825 65.36 0.96 ;
        RECT 65.2875 0.315 65.3575 0.9625 ;
        RECT 64.835 0.315 65.3575 0.385 ;
        RECT 64.835 0.2825 64.905 0.4175 ;
      LAYER via1 ;
        RECT 64.8375 0.3175 64.9025 0.3825 ;
        RECT 65.2925 0.86 65.3575 0.925 ;
      LAYER via2 ;
        RECT 65.2875 0.8575 65.3575 0.9275 ;
    END
  END rs2_sel[18]
  PIN rs2_sel[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 68.7525 0.8225 68.8225 0.9625 ;
      LAYER metal1 ;
        RECT 68.7575 0.825 68.8225 0.96 ;
        RECT 68.3025 0.2825 68.3675 0.4175 ;
      LAYER metal2 ;
        RECT 68.7525 0.825 68.825 0.96 ;
        RECT 68.7525 0.315 68.8225 0.9625 ;
        RECT 68.3 0.315 68.8225 0.385 ;
        RECT 68.3 0.2825 68.37 0.4175 ;
      LAYER via1 ;
        RECT 68.3025 0.3175 68.3675 0.3825 ;
        RECT 68.7575 0.86 68.8225 0.925 ;
      LAYER via2 ;
        RECT 68.7525 0.8575 68.8225 0.9275 ;
    END
  END rs2_sel[19]
  PIN rs2_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 6.3825 0.8225 6.4525 0.9625 ;
      LAYER metal1 ;
        RECT 6.3875 0.825 6.4525 0.96 ;
        RECT 5.9325 0.2825 5.9975 0.4175 ;
      LAYER metal2 ;
        RECT 6.3825 0.825 6.455 0.96 ;
        RECT 6.3825 0.315 6.4525 0.9625 ;
        RECT 5.93 0.315 6.4525 0.385 ;
        RECT 5.93 0.2825 6 0.4175 ;
      LAYER via1 ;
        RECT 5.9325 0.3175 5.9975 0.3825 ;
        RECT 6.3875 0.86 6.4525 0.925 ;
      LAYER via2 ;
        RECT 6.3825 0.8575 6.4525 0.9275 ;
    END
  END rs2_sel[1]
  PIN rs2_sel[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 72.2175 0.8225 72.2875 0.9625 ;
      LAYER metal1 ;
        RECT 72.2225 0.825 72.2875 0.96 ;
        RECT 71.7675 0.2825 71.8325 0.4175 ;
      LAYER metal2 ;
        RECT 72.2175 0.825 72.29 0.96 ;
        RECT 72.2175 0.315 72.2875 0.9625 ;
        RECT 71.765 0.315 72.2875 0.385 ;
        RECT 71.765 0.2825 71.835 0.4175 ;
      LAYER via1 ;
        RECT 71.7675 0.3175 71.8325 0.3825 ;
        RECT 72.2225 0.86 72.2875 0.925 ;
      LAYER via2 ;
        RECT 72.2175 0.8575 72.2875 0.9275 ;
    END
  END rs2_sel[20]
  PIN rs2_sel[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.6825 0.8225 75.7525 0.9625 ;
      LAYER metal1 ;
        RECT 75.6875 0.825 75.7525 0.96 ;
        RECT 75.2325 0.2825 75.2975 0.4175 ;
      LAYER metal2 ;
        RECT 75.6825 0.825 75.755 0.96 ;
        RECT 75.6825 0.315 75.7525 0.9625 ;
        RECT 75.23 0.315 75.7525 0.385 ;
        RECT 75.23 0.2825 75.3 0.4175 ;
      LAYER via1 ;
        RECT 75.2325 0.3175 75.2975 0.3825 ;
        RECT 75.6875 0.86 75.7525 0.925 ;
      LAYER via2 ;
        RECT 75.6825 0.8575 75.7525 0.9275 ;
    END
  END rs2_sel[21]
  PIN rs2_sel[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 79.1475 0.8225 79.2175 0.9625 ;
      LAYER metal1 ;
        RECT 79.1525 0.825 79.2175 0.96 ;
        RECT 78.6975 0.2825 78.7625 0.4175 ;
      LAYER metal2 ;
        RECT 79.1475 0.825 79.22 0.96 ;
        RECT 79.1475 0.315 79.2175 0.9625 ;
        RECT 78.695 0.315 79.2175 0.385 ;
        RECT 78.695 0.2825 78.765 0.4175 ;
      LAYER via1 ;
        RECT 78.6975 0.3175 78.7625 0.3825 ;
        RECT 79.1525 0.86 79.2175 0.925 ;
      LAYER via2 ;
        RECT 79.1475 0.8575 79.2175 0.9275 ;
    END
  END rs2_sel[22]
  PIN rs2_sel[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 82.6125 0.8225 82.6825 0.9625 ;
      LAYER metal1 ;
        RECT 82.6175 0.825 82.6825 0.96 ;
        RECT 82.1625 0.2825 82.2275 0.4175 ;
      LAYER metal2 ;
        RECT 82.6125 0.825 82.685 0.96 ;
        RECT 82.6125 0.315 82.6825 0.9625 ;
        RECT 82.16 0.315 82.6825 0.385 ;
        RECT 82.16 0.2825 82.23 0.4175 ;
      LAYER via1 ;
        RECT 82.1625 0.3175 82.2275 0.3825 ;
        RECT 82.6175 0.86 82.6825 0.925 ;
      LAYER via2 ;
        RECT 82.6125 0.8575 82.6825 0.9275 ;
    END
  END rs2_sel[23]
  PIN rs2_sel[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 86.0775 0.8225 86.1475 0.9625 ;
      LAYER metal1 ;
        RECT 86.0825 0.825 86.1475 0.96 ;
        RECT 85.6275 0.2825 85.6925 0.4175 ;
      LAYER metal2 ;
        RECT 86.0775 0.825 86.15 0.96 ;
        RECT 86.0775 0.315 86.1475 0.9625 ;
        RECT 85.625 0.315 86.1475 0.385 ;
        RECT 85.625 0.2825 85.695 0.4175 ;
      LAYER via1 ;
        RECT 85.6275 0.3175 85.6925 0.3825 ;
        RECT 86.0825 0.86 86.1475 0.925 ;
      LAYER via2 ;
        RECT 86.0775 0.8575 86.1475 0.9275 ;
    END
  END rs2_sel[24]
  PIN rs2_sel[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 89.5425 0.8225 89.6125 0.9625 ;
      LAYER metal1 ;
        RECT 89.5475 0.825 89.6125 0.96 ;
        RECT 89.0925 0.2825 89.1575 0.4175 ;
      LAYER metal2 ;
        RECT 89.5425 0.825 89.615 0.96 ;
        RECT 89.5425 0.315 89.6125 0.9625 ;
        RECT 89.09 0.315 89.6125 0.385 ;
        RECT 89.09 0.2825 89.16 0.4175 ;
      LAYER via1 ;
        RECT 89.0925 0.3175 89.1575 0.3825 ;
        RECT 89.5475 0.86 89.6125 0.925 ;
      LAYER via2 ;
        RECT 89.5425 0.8575 89.6125 0.9275 ;
    END
  END rs2_sel[25]
  PIN rs2_sel[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 93.0075 0.8225 93.0775 0.9625 ;
      LAYER metal1 ;
        RECT 93.0125 0.825 93.0775 0.96 ;
        RECT 92.5575 0.2825 92.6225 0.4175 ;
      LAYER metal2 ;
        RECT 93.0075 0.825 93.08 0.96 ;
        RECT 93.0075 0.315 93.0775 0.9625 ;
        RECT 92.555 0.315 93.0775 0.385 ;
        RECT 92.555 0.2825 92.625 0.4175 ;
      LAYER via1 ;
        RECT 92.5575 0.3175 92.6225 0.3825 ;
        RECT 93.0125 0.86 93.0775 0.925 ;
      LAYER via2 ;
        RECT 93.0075 0.8575 93.0775 0.9275 ;
    END
  END rs2_sel[26]
  PIN rs2_sel[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 96.4725 0.8225 96.5425 0.9625 ;
      LAYER metal1 ;
        RECT 96.4775 0.825 96.5425 0.96 ;
        RECT 96.0225 0.2825 96.0875 0.4175 ;
      LAYER metal2 ;
        RECT 96.4725 0.825 96.545 0.96 ;
        RECT 96.4725 0.315 96.5425 0.9625 ;
        RECT 96.02 0.315 96.5425 0.385 ;
        RECT 96.02 0.2825 96.09 0.4175 ;
      LAYER via1 ;
        RECT 96.0225 0.3175 96.0875 0.3825 ;
        RECT 96.4775 0.86 96.5425 0.925 ;
      LAYER via2 ;
        RECT 96.4725 0.8575 96.5425 0.9275 ;
    END
  END rs2_sel[27]
  PIN rs2_sel[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 99.9375 0.8225 100.0075 0.9625 ;
      LAYER metal1 ;
        RECT 99.9425 0.825 100.0075 0.96 ;
        RECT 99.4875 0.2825 99.5525 0.4175 ;
      LAYER metal2 ;
        RECT 99.9375 0.825 100.01 0.96 ;
        RECT 99.9375 0.315 100.0075 0.9625 ;
        RECT 99.485 0.315 100.0075 0.385 ;
        RECT 99.485 0.2825 99.555 0.4175 ;
      LAYER via1 ;
        RECT 99.4875 0.3175 99.5525 0.3825 ;
        RECT 99.9425 0.86 100.0075 0.925 ;
      LAYER via2 ;
        RECT 99.9375 0.8575 100.0075 0.9275 ;
    END
  END rs2_sel[28]
  PIN rs2_sel[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 103.4025 0.8225 103.4725 0.9625 ;
      LAYER metal1 ;
        RECT 103.4075 0.825 103.4725 0.96 ;
        RECT 102.9525 0.2825 103.0175 0.4175 ;
      LAYER metal2 ;
        RECT 103.4025 0.825 103.475 0.96 ;
        RECT 103.4025 0.315 103.4725 0.9625 ;
        RECT 102.95 0.315 103.4725 0.385 ;
        RECT 102.95 0.2825 103.02 0.4175 ;
      LAYER via1 ;
        RECT 102.9525 0.3175 103.0175 0.3825 ;
        RECT 103.4075 0.86 103.4725 0.925 ;
      LAYER via2 ;
        RECT 103.4025 0.8575 103.4725 0.9275 ;
    END
  END rs2_sel[29]
  PIN rs2_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 9.8475 0.8225 9.9175 0.9625 ;
      LAYER metal1 ;
        RECT 9.8525 0.825 9.9175 0.96 ;
        RECT 9.3975 0.2825 9.4625 0.4175 ;
      LAYER metal2 ;
        RECT 9.8475 0.825 9.92 0.96 ;
        RECT 9.8475 0.315 9.9175 0.9625 ;
        RECT 9.395 0.315 9.9175 0.385 ;
        RECT 9.395 0.2825 9.465 0.4175 ;
      LAYER via1 ;
        RECT 9.3975 0.3175 9.4625 0.3825 ;
        RECT 9.8525 0.86 9.9175 0.925 ;
      LAYER via2 ;
        RECT 9.8475 0.8575 9.9175 0.9275 ;
    END
  END rs2_sel[2]
  PIN rs2_sel[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 106.8675 0.8225 106.9375 0.9625 ;
      LAYER metal1 ;
        RECT 106.8725 0.825 106.9375 0.96 ;
        RECT 106.4175 0.2825 106.4825 0.4175 ;
      LAYER metal2 ;
        RECT 106.8675 0.825 106.94 0.96 ;
        RECT 106.8675 0.315 106.9375 0.9625 ;
        RECT 106.415 0.315 106.9375 0.385 ;
        RECT 106.415 0.2825 106.485 0.4175 ;
      LAYER via1 ;
        RECT 106.4175 0.3175 106.4825 0.3825 ;
        RECT 106.8725 0.86 106.9375 0.925 ;
      LAYER via2 ;
        RECT 106.8675 0.8575 106.9375 0.9275 ;
    END
  END rs2_sel[30]
  PIN rs2_sel[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 110.3325 0.8225 110.4025 0.9625 ;
      LAYER metal1 ;
        RECT 110.3375 0.825 110.4025 0.96 ;
        RECT 109.8825 0.2825 109.9475 0.4175 ;
      LAYER metal2 ;
        RECT 110.3325 0.825 110.405 0.96 ;
        RECT 110.3325 0.315 110.4025 0.9625 ;
        RECT 109.88 0.315 110.4025 0.385 ;
        RECT 109.88 0.2825 109.95 0.4175 ;
      LAYER via1 ;
        RECT 109.8825 0.3175 109.9475 0.3825 ;
        RECT 110.3375 0.86 110.4025 0.925 ;
      LAYER via2 ;
        RECT 110.3325 0.8575 110.4025 0.9275 ;
    END
  END rs2_sel[31]
  PIN rs2_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 13.3125 0.8225 13.3825 0.9625 ;
      LAYER metal1 ;
        RECT 13.3175 0.825 13.3825 0.96 ;
        RECT 12.8625 0.2825 12.9275 0.4175 ;
      LAYER metal2 ;
        RECT 13.3125 0.825 13.385 0.96 ;
        RECT 13.3125 0.315 13.3825 0.9625 ;
        RECT 12.86 0.315 13.3825 0.385 ;
        RECT 12.86 0.2825 12.93 0.4175 ;
      LAYER via1 ;
        RECT 12.8625 0.3175 12.9275 0.3825 ;
        RECT 13.3175 0.86 13.3825 0.925 ;
      LAYER via2 ;
        RECT 13.3125 0.8575 13.3825 0.9275 ;
    END
  END rs2_sel[3]
  PIN rs2_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 16.7775 0.8225 16.8475 0.9625 ;
      LAYER metal1 ;
        RECT 16.7825 0.825 16.8475 0.96 ;
        RECT 16.3275 0.2825 16.3925 0.4175 ;
      LAYER metal2 ;
        RECT 16.7775 0.825 16.85 0.96 ;
        RECT 16.7775 0.315 16.8475 0.9625 ;
        RECT 16.325 0.315 16.8475 0.385 ;
        RECT 16.325 0.2825 16.395 0.4175 ;
      LAYER via1 ;
        RECT 16.3275 0.3175 16.3925 0.3825 ;
        RECT 16.7825 0.86 16.8475 0.925 ;
      LAYER via2 ;
        RECT 16.7775 0.8575 16.8475 0.9275 ;
    END
  END rs2_sel[4]
  PIN rs2_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 20.2425 0.8225 20.3125 0.9625 ;
      LAYER metal1 ;
        RECT 20.2475 0.825 20.3125 0.96 ;
        RECT 19.7925 0.2825 19.8575 0.4175 ;
      LAYER metal2 ;
        RECT 20.2425 0.825 20.315 0.96 ;
        RECT 20.2425 0.315 20.3125 0.9625 ;
        RECT 19.79 0.315 20.3125 0.385 ;
        RECT 19.79 0.2825 19.86 0.4175 ;
      LAYER via1 ;
        RECT 19.7925 0.3175 19.8575 0.3825 ;
        RECT 20.2475 0.86 20.3125 0.925 ;
      LAYER via2 ;
        RECT 20.2425 0.8575 20.3125 0.9275 ;
    END
  END rs2_sel[5]
  PIN rs2_sel[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 23.7075 0.8225 23.7775 0.9625 ;
      LAYER metal1 ;
        RECT 23.7125 0.825 23.7775 0.96 ;
        RECT 23.2575 0.2825 23.3225 0.4175 ;
      LAYER metal2 ;
        RECT 23.7075 0.825 23.78 0.96 ;
        RECT 23.7075 0.315 23.7775 0.9625 ;
        RECT 23.255 0.315 23.7775 0.385 ;
        RECT 23.255 0.2825 23.325 0.4175 ;
      LAYER via1 ;
        RECT 23.2575 0.3175 23.3225 0.3825 ;
        RECT 23.7125 0.86 23.7775 0.925 ;
      LAYER via2 ;
        RECT 23.7075 0.8575 23.7775 0.9275 ;
    END
  END rs2_sel[6]
  PIN rs2_sel[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 27.1725 0.8225 27.2425 0.9625 ;
      LAYER metal1 ;
        RECT 27.1775 0.825 27.2425 0.96 ;
        RECT 26.7225 0.2825 26.7875 0.4175 ;
      LAYER metal2 ;
        RECT 27.1725 0.825 27.245 0.96 ;
        RECT 27.1725 0.315 27.2425 0.9625 ;
        RECT 26.72 0.315 27.2425 0.385 ;
        RECT 26.72 0.2825 26.79 0.4175 ;
      LAYER via1 ;
        RECT 26.7225 0.3175 26.7875 0.3825 ;
        RECT 27.1775 0.86 27.2425 0.925 ;
      LAYER via2 ;
        RECT 27.1725 0.8575 27.2425 0.9275 ;
    END
  END rs2_sel[7]
  PIN rs2_sel[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 30.6375 0.8225 30.7075 0.9625 ;
      LAYER metal1 ;
        RECT 30.6425 0.825 30.7075 0.96 ;
        RECT 30.1875 0.2825 30.2525 0.4175 ;
      LAYER metal2 ;
        RECT 30.6375 0.825 30.71 0.96 ;
        RECT 30.6375 0.315 30.7075 0.9625 ;
        RECT 30.185 0.315 30.7075 0.385 ;
        RECT 30.185 0.2825 30.255 0.4175 ;
      LAYER via1 ;
        RECT 30.1875 0.3175 30.2525 0.3825 ;
        RECT 30.6425 0.86 30.7075 0.925 ;
      LAYER via2 ;
        RECT 30.6375 0.8575 30.7075 0.9275 ;
    END
  END rs2_sel[8]
  PIN rs2_sel[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 34.1025 0.8225 34.1725 0.9625 ;
      LAYER metal1 ;
        RECT 34.1075 0.825 34.1725 0.96 ;
        RECT 33.6525 0.2825 33.7175 0.4175 ;
      LAYER metal2 ;
        RECT 34.1025 0.825 34.175 0.96 ;
        RECT 34.1025 0.315 34.1725 0.9625 ;
        RECT 33.65 0.315 34.1725 0.385 ;
        RECT 33.65 0.2825 33.72 0.4175 ;
      LAYER via1 ;
        RECT 33.6525 0.3175 33.7175 0.3825 ;
        RECT 34.1075 0.86 34.1725 0.925 ;
      LAYER via2 ;
        RECT 34.1025 0.8575 34.1725 0.9275 ;
    END
  END rs2_sel[9]
  OBS
    LAYER metal1 ;
      RECT 114.3225 1.22 114.3875 1.355 ;
      RECT 114.32 0.265 114.385 1.3325 ;
      RECT 114.32 0.265 114.3875 0.4 ;
      RECT 113.6025 1.2075 113.67 1.3425 ;
      RECT 113.605 0.265 113.67 1.3425 ;
      RECT 113.6025 0.265 113.67 0.4 ;
      RECT 113.415 1.2075 113.4825 1.3425 ;
      RECT 113.415 0.265 113.48 1.3425 ;
      RECT 113.415 0.265 113.4825 0.4 ;
      RECT 112.6975 1.22 112.7625 1.355 ;
      RECT 112.7 0.265 112.765 1.3325 ;
      RECT 112.6975 0.265 112.765 0.4 ;
      RECT 111.515 0.265 111.58 1.3725 ;
      RECT 111.515 0.4625 111.6025 0.5975 ;
      RECT 111.13 0.28 111.195 1.3725 ;
      RECT 111.13 0.72 111.2175 0.855 ;
      RECT 110.565 0.265 110.63 1.3725 ;
      RECT 110.5425 0.725 110.63 0.86 ;
      RECT 110.1575 1.2375 110.245 1.3725 ;
      RECT 110.18 0.28 110.245 1.3725 ;
      RECT 109.975 0.4875 110.04 1.14 ;
      RECT 109.975 0.6825 110.0725 0.8175 ;
      RECT 109.785 0.4875 109.85 1.14 ;
      RECT 109.7675 0.8675 109.85 1.0025 ;
      RECT 109.6 0.4875 109.665 1.14 ;
      RECT 109.6 0.8675 109.6825 1.0025 ;
      RECT 109.41 0.485 109.475 1.14 ;
      RECT 109.3775 0.4675 109.4425 0.6025 ;
      RECT 109.025 0.28 109.09 1.3725 ;
      RECT 109.0025 0.6625 109.09 0.7975 ;
      RECT 108.82 0.28 108.885 1.3725 ;
      RECT 108.82 0.8675 108.9075 1.0025 ;
      RECT 108.445 0.4875 108.51 1.14 ;
      RECT 108.445 0.6625 108.5275 0.7975 ;
      RECT 108.255 0.4875 108.32 1.14 ;
      RECT 108.2225 0.87 108.32 1.005 ;
      RECT 108.05 0.4875 108.115 1.14 ;
      RECT 108.05 0.87 108.1475 1.005 ;
      RECT 107.6875 1.25 107.7525 1.385 ;
      RECT 107.665 0.28 107.73 1.3725 ;
      RECT 107.1 0.265 107.165 1.3725 ;
      RECT 107.0775 0.725 107.165 0.86 ;
      RECT 106.6925 1.2375 106.78 1.3725 ;
      RECT 106.715 0.28 106.78 1.3725 ;
      RECT 106.51 0.4875 106.575 1.14 ;
      RECT 106.51 0.6825 106.6075 0.8175 ;
      RECT 106.32 0.4875 106.385 1.14 ;
      RECT 106.3025 0.8675 106.385 1.0025 ;
      RECT 106.135 0.4875 106.2 1.14 ;
      RECT 106.135 0.8675 106.2175 1.0025 ;
      RECT 105.945 0.485 106.01 1.14 ;
      RECT 105.9125 0.4675 105.9775 0.6025 ;
      RECT 105.56 0.28 105.625 1.3725 ;
      RECT 105.5375 0.6625 105.625 0.7975 ;
      RECT 105.355 0.28 105.42 1.3725 ;
      RECT 105.355 0.8675 105.4425 1.0025 ;
      RECT 104.98 0.4875 105.045 1.14 ;
      RECT 104.98 0.6625 105.0625 0.7975 ;
      RECT 104.79 0.4875 104.855 1.14 ;
      RECT 104.7575 0.87 104.855 1.005 ;
      RECT 104.585 0.4875 104.65 1.14 ;
      RECT 104.585 0.87 104.6825 1.005 ;
      RECT 104.2225 1.25 104.2875 1.385 ;
      RECT 104.2 0.28 104.265 1.3725 ;
      RECT 103.635 0.265 103.7 1.3725 ;
      RECT 103.6125 0.725 103.7 0.86 ;
      RECT 103.2275 1.2375 103.315 1.3725 ;
      RECT 103.25 0.28 103.315 1.3725 ;
      RECT 103.045 0.4875 103.11 1.14 ;
      RECT 103.045 0.6825 103.1425 0.8175 ;
      RECT 102.855 0.4875 102.92 1.14 ;
      RECT 102.8375 0.8675 102.92 1.0025 ;
      RECT 102.67 0.4875 102.735 1.14 ;
      RECT 102.67 0.8675 102.7525 1.0025 ;
      RECT 102.48 0.485 102.545 1.14 ;
      RECT 102.4475 0.4675 102.5125 0.6025 ;
      RECT 102.095 0.28 102.16 1.3725 ;
      RECT 102.0725 0.6625 102.16 0.7975 ;
      RECT 101.89 0.28 101.955 1.3725 ;
      RECT 101.89 0.8675 101.9775 1.0025 ;
      RECT 101.515 0.4875 101.58 1.14 ;
      RECT 101.515 0.6625 101.5975 0.7975 ;
      RECT 101.325 0.4875 101.39 1.14 ;
      RECT 101.2925 0.87 101.39 1.005 ;
      RECT 101.12 0.4875 101.185 1.14 ;
      RECT 101.12 0.87 101.2175 1.005 ;
      RECT 100.7575 1.25 100.8225 1.385 ;
      RECT 100.735 0.28 100.8 1.3725 ;
      RECT 100.17 0.265 100.235 1.3725 ;
      RECT 100.1475 0.725 100.235 0.86 ;
      RECT 99.7625 1.2375 99.85 1.3725 ;
      RECT 99.785 0.28 99.85 1.3725 ;
      RECT 99.58 0.4875 99.645 1.14 ;
      RECT 99.58 0.6825 99.6775 0.8175 ;
      RECT 99.39 0.4875 99.455 1.14 ;
      RECT 99.3725 0.8675 99.455 1.0025 ;
      RECT 99.205 0.4875 99.27 1.14 ;
      RECT 99.205 0.8675 99.2875 1.0025 ;
      RECT 99.015 0.485 99.08 1.14 ;
      RECT 98.9825 0.4675 99.0475 0.6025 ;
      RECT 98.63 0.28 98.695 1.3725 ;
      RECT 98.6075 0.6625 98.695 0.7975 ;
      RECT 98.425 0.28 98.49 1.3725 ;
      RECT 98.425 0.8675 98.5125 1.0025 ;
      RECT 98.05 0.4875 98.115 1.14 ;
      RECT 98.05 0.6625 98.1325 0.7975 ;
      RECT 97.86 0.4875 97.925 1.14 ;
      RECT 97.8275 0.87 97.925 1.005 ;
      RECT 97.655 0.4875 97.72 1.14 ;
      RECT 97.655 0.87 97.7525 1.005 ;
      RECT 97.2925 1.25 97.3575 1.385 ;
      RECT 97.27 0.28 97.335 1.3725 ;
      RECT 96.705 0.265 96.77 1.3725 ;
      RECT 96.6825 0.725 96.77 0.86 ;
      RECT 96.2975 1.2375 96.385 1.3725 ;
      RECT 96.32 0.28 96.385 1.3725 ;
      RECT 96.115 0.4875 96.18 1.14 ;
      RECT 96.115 0.6825 96.2125 0.8175 ;
      RECT 95.925 0.4875 95.99 1.14 ;
      RECT 95.9075 0.8675 95.99 1.0025 ;
      RECT 95.74 0.4875 95.805 1.14 ;
      RECT 95.74 0.8675 95.8225 1.0025 ;
      RECT 95.55 0.485 95.615 1.14 ;
      RECT 95.5175 0.4675 95.5825 0.6025 ;
      RECT 95.165 0.28 95.23 1.3725 ;
      RECT 95.1425 0.6625 95.23 0.7975 ;
      RECT 94.96 0.28 95.025 1.3725 ;
      RECT 94.96 0.8675 95.0475 1.0025 ;
      RECT 94.585 0.4875 94.65 1.14 ;
      RECT 94.585 0.6625 94.6675 0.7975 ;
      RECT 94.395 0.4875 94.46 1.14 ;
      RECT 94.3625 0.87 94.46 1.005 ;
      RECT 94.19 0.4875 94.255 1.14 ;
      RECT 94.19 0.87 94.2875 1.005 ;
      RECT 93.8275 1.25 93.8925 1.385 ;
      RECT 93.805 0.28 93.87 1.3725 ;
      RECT 93.24 0.265 93.305 1.3725 ;
      RECT 93.2175 0.725 93.305 0.86 ;
      RECT 92.8325 1.2375 92.92 1.3725 ;
      RECT 92.855 0.28 92.92 1.3725 ;
      RECT 92.65 0.4875 92.715 1.14 ;
      RECT 92.65 0.6825 92.7475 0.8175 ;
      RECT 92.46 0.4875 92.525 1.14 ;
      RECT 92.4425 0.8675 92.525 1.0025 ;
      RECT 92.275 0.4875 92.34 1.14 ;
      RECT 92.275 0.8675 92.3575 1.0025 ;
      RECT 92.085 0.485 92.15 1.14 ;
      RECT 92.0525 0.4675 92.1175 0.6025 ;
      RECT 91.7 0.28 91.765 1.3725 ;
      RECT 91.6775 0.6625 91.765 0.7975 ;
      RECT 91.495 0.28 91.56 1.3725 ;
      RECT 91.495 0.8675 91.5825 1.0025 ;
      RECT 91.12 0.4875 91.185 1.14 ;
      RECT 91.12 0.6625 91.2025 0.7975 ;
      RECT 90.93 0.4875 90.995 1.14 ;
      RECT 90.8975 0.87 90.995 1.005 ;
      RECT 90.725 0.4875 90.79 1.14 ;
      RECT 90.725 0.87 90.8225 1.005 ;
      RECT 90.3625 1.25 90.4275 1.385 ;
      RECT 90.34 0.28 90.405 1.3725 ;
      RECT 89.775 0.265 89.84 1.3725 ;
      RECT 89.7525 0.725 89.84 0.86 ;
      RECT 89.3675 1.2375 89.455 1.3725 ;
      RECT 89.39 0.28 89.455 1.3725 ;
      RECT 89.185 0.4875 89.25 1.14 ;
      RECT 89.185 0.6825 89.2825 0.8175 ;
      RECT 88.995 0.4875 89.06 1.14 ;
      RECT 88.9775 0.8675 89.06 1.0025 ;
      RECT 88.81 0.4875 88.875 1.14 ;
      RECT 88.81 0.8675 88.8925 1.0025 ;
      RECT 88.62 0.485 88.685 1.14 ;
      RECT 88.5875 0.4675 88.6525 0.6025 ;
      RECT 88.235 0.28 88.3 1.3725 ;
      RECT 88.2125 0.6625 88.3 0.7975 ;
      RECT 88.03 0.28 88.095 1.3725 ;
      RECT 88.03 0.8675 88.1175 1.0025 ;
      RECT 87.655 0.4875 87.72 1.14 ;
      RECT 87.655 0.6625 87.7375 0.7975 ;
      RECT 87.465 0.4875 87.53 1.14 ;
      RECT 87.4325 0.87 87.53 1.005 ;
      RECT 87.26 0.4875 87.325 1.14 ;
      RECT 87.26 0.87 87.3575 1.005 ;
      RECT 86.8975 1.25 86.9625 1.385 ;
      RECT 86.875 0.28 86.94 1.3725 ;
      RECT 86.31 0.265 86.375 1.3725 ;
      RECT 86.2875 0.725 86.375 0.86 ;
      RECT 85.9025 1.2375 85.99 1.3725 ;
      RECT 85.925 0.28 85.99 1.3725 ;
      RECT 85.72 0.4875 85.785 1.14 ;
      RECT 85.72 0.6825 85.8175 0.8175 ;
      RECT 85.53 0.4875 85.595 1.14 ;
      RECT 85.5125 0.8675 85.595 1.0025 ;
      RECT 85.345 0.4875 85.41 1.14 ;
      RECT 85.345 0.8675 85.4275 1.0025 ;
      RECT 85.155 0.485 85.22 1.14 ;
      RECT 85.1225 0.4675 85.1875 0.6025 ;
      RECT 84.77 0.28 84.835 1.3725 ;
      RECT 84.7475 0.6625 84.835 0.7975 ;
      RECT 84.565 0.28 84.63 1.3725 ;
      RECT 84.565 0.8675 84.6525 1.0025 ;
      RECT 84.19 0.4875 84.255 1.14 ;
      RECT 84.19 0.6625 84.2725 0.7975 ;
      RECT 84 0.4875 84.065 1.14 ;
      RECT 83.9675 0.87 84.065 1.005 ;
      RECT 83.795 0.4875 83.86 1.14 ;
      RECT 83.795 0.87 83.8925 1.005 ;
      RECT 83.4325 1.25 83.4975 1.385 ;
      RECT 83.41 0.28 83.475 1.3725 ;
      RECT 82.845 0.265 82.91 1.3725 ;
      RECT 82.8225 0.725 82.91 0.86 ;
      RECT 82.4375 1.2375 82.525 1.3725 ;
      RECT 82.46 0.28 82.525 1.3725 ;
      RECT 82.255 0.4875 82.32 1.14 ;
      RECT 82.255 0.6825 82.3525 0.8175 ;
      RECT 82.065 0.4875 82.13 1.14 ;
      RECT 82.0475 0.8675 82.13 1.0025 ;
      RECT 81.88 0.4875 81.945 1.14 ;
      RECT 81.88 0.8675 81.9625 1.0025 ;
      RECT 81.69 0.485 81.755 1.14 ;
      RECT 81.6575 0.4675 81.7225 0.6025 ;
      RECT 81.305 0.28 81.37 1.3725 ;
      RECT 81.2825 0.6625 81.37 0.7975 ;
      RECT 81.1 0.28 81.165 1.3725 ;
      RECT 81.1 0.8675 81.1875 1.0025 ;
      RECT 80.725 0.4875 80.79 1.14 ;
      RECT 80.725 0.6625 80.8075 0.7975 ;
      RECT 80.535 0.4875 80.6 1.14 ;
      RECT 80.5025 0.87 80.6 1.005 ;
      RECT 80.33 0.4875 80.395 1.14 ;
      RECT 80.33 0.87 80.4275 1.005 ;
      RECT 79.9675 1.25 80.0325 1.385 ;
      RECT 79.945 0.28 80.01 1.3725 ;
      RECT 79.38 0.265 79.445 1.3725 ;
      RECT 79.3575 0.725 79.445 0.86 ;
      RECT 78.9725 1.2375 79.06 1.3725 ;
      RECT 78.995 0.28 79.06 1.3725 ;
      RECT 78.79 0.4875 78.855 1.14 ;
      RECT 78.79 0.6825 78.8875 0.8175 ;
      RECT 78.6 0.4875 78.665 1.14 ;
      RECT 78.5825 0.8675 78.665 1.0025 ;
      RECT 78.415 0.4875 78.48 1.14 ;
      RECT 78.415 0.8675 78.4975 1.0025 ;
      RECT 78.225 0.485 78.29 1.14 ;
      RECT 78.1925 0.4675 78.2575 0.6025 ;
      RECT 77.84 0.28 77.905 1.3725 ;
      RECT 77.8175 0.6625 77.905 0.7975 ;
      RECT 77.635 0.28 77.7 1.3725 ;
      RECT 77.635 0.8675 77.7225 1.0025 ;
      RECT 77.26 0.4875 77.325 1.14 ;
      RECT 77.26 0.6625 77.3425 0.7975 ;
      RECT 77.07 0.4875 77.135 1.14 ;
      RECT 77.0375 0.87 77.135 1.005 ;
      RECT 76.865 0.4875 76.93 1.14 ;
      RECT 76.865 0.87 76.9625 1.005 ;
      RECT 76.5025 1.25 76.5675 1.385 ;
      RECT 76.48 0.28 76.545 1.3725 ;
      RECT 75.915 0.265 75.98 1.3725 ;
      RECT 75.8925 0.725 75.98 0.86 ;
      RECT 75.5075 1.2375 75.595 1.3725 ;
      RECT 75.53 0.28 75.595 1.3725 ;
      RECT 75.325 0.4875 75.39 1.14 ;
      RECT 75.325 0.6825 75.4225 0.8175 ;
      RECT 75.135 0.4875 75.2 1.14 ;
      RECT 75.1175 0.8675 75.2 1.0025 ;
      RECT 74.95 0.4875 75.015 1.14 ;
      RECT 74.95 0.8675 75.0325 1.0025 ;
      RECT 74.76 0.485 74.825 1.14 ;
      RECT 74.7275 0.4675 74.7925 0.6025 ;
      RECT 74.375 0.28 74.44 1.3725 ;
      RECT 74.3525 0.6625 74.44 0.7975 ;
      RECT 74.17 0.28 74.235 1.3725 ;
      RECT 74.17 0.8675 74.2575 1.0025 ;
      RECT 73.795 0.4875 73.86 1.14 ;
      RECT 73.795 0.6625 73.8775 0.7975 ;
      RECT 73.605 0.4875 73.67 1.14 ;
      RECT 73.5725 0.87 73.67 1.005 ;
      RECT 73.4 0.4875 73.465 1.14 ;
      RECT 73.4 0.87 73.4975 1.005 ;
      RECT 73.0375 1.25 73.1025 1.385 ;
      RECT 73.015 0.28 73.08 1.3725 ;
      RECT 72.45 0.265 72.515 1.3725 ;
      RECT 72.4275 0.725 72.515 0.86 ;
      RECT 72.0425 1.2375 72.13 1.3725 ;
      RECT 72.065 0.28 72.13 1.3725 ;
      RECT 71.86 0.4875 71.925 1.14 ;
      RECT 71.86 0.6825 71.9575 0.8175 ;
      RECT 71.67 0.4875 71.735 1.14 ;
      RECT 71.6525 0.8675 71.735 1.0025 ;
      RECT 71.485 0.4875 71.55 1.14 ;
      RECT 71.485 0.8675 71.5675 1.0025 ;
      RECT 71.295 0.485 71.36 1.14 ;
      RECT 71.2625 0.4675 71.3275 0.6025 ;
      RECT 70.91 0.28 70.975 1.3725 ;
      RECT 70.8875 0.6625 70.975 0.7975 ;
      RECT 70.705 0.28 70.77 1.3725 ;
      RECT 70.705 0.8675 70.7925 1.0025 ;
      RECT 70.33 0.4875 70.395 1.14 ;
      RECT 70.33 0.6625 70.4125 0.7975 ;
      RECT 70.14 0.4875 70.205 1.14 ;
      RECT 70.1075 0.87 70.205 1.005 ;
      RECT 69.935 0.4875 70 1.14 ;
      RECT 69.935 0.87 70.0325 1.005 ;
      RECT 69.5725 1.25 69.6375 1.385 ;
      RECT 69.55 0.28 69.615 1.3725 ;
      RECT 68.985 0.265 69.05 1.3725 ;
      RECT 68.9625 0.725 69.05 0.86 ;
      RECT 68.5775 1.2375 68.665 1.3725 ;
      RECT 68.6 0.28 68.665 1.3725 ;
      RECT 68.395 0.4875 68.46 1.14 ;
      RECT 68.395 0.6825 68.4925 0.8175 ;
      RECT 68.205 0.4875 68.27 1.14 ;
      RECT 68.1875 0.8675 68.27 1.0025 ;
      RECT 68.02 0.4875 68.085 1.14 ;
      RECT 68.02 0.8675 68.1025 1.0025 ;
      RECT 67.83 0.485 67.895 1.14 ;
      RECT 67.7975 0.4675 67.8625 0.6025 ;
      RECT 67.445 0.28 67.51 1.3725 ;
      RECT 67.4225 0.6625 67.51 0.7975 ;
      RECT 67.24 0.28 67.305 1.3725 ;
      RECT 67.24 0.8675 67.3275 1.0025 ;
      RECT 66.865 0.4875 66.93 1.14 ;
      RECT 66.865 0.6625 66.9475 0.7975 ;
      RECT 66.675 0.4875 66.74 1.14 ;
      RECT 66.6425 0.87 66.74 1.005 ;
      RECT 66.47 0.4875 66.535 1.14 ;
      RECT 66.47 0.87 66.5675 1.005 ;
      RECT 66.1075 1.25 66.1725 1.385 ;
      RECT 66.085 0.28 66.15 1.3725 ;
      RECT 65.52 0.265 65.585 1.3725 ;
      RECT 65.4975 0.725 65.585 0.86 ;
      RECT 65.1125 1.2375 65.2 1.3725 ;
      RECT 65.135 0.28 65.2 1.3725 ;
      RECT 64.93 0.4875 64.995 1.14 ;
      RECT 64.93 0.6825 65.0275 0.8175 ;
      RECT 64.74 0.4875 64.805 1.14 ;
      RECT 64.7225 0.8675 64.805 1.0025 ;
      RECT 64.555 0.4875 64.62 1.14 ;
      RECT 64.555 0.8675 64.6375 1.0025 ;
      RECT 64.365 0.485 64.43 1.14 ;
      RECT 64.3325 0.4675 64.3975 0.6025 ;
      RECT 63.98 0.28 64.045 1.3725 ;
      RECT 63.9575 0.6625 64.045 0.7975 ;
      RECT 63.775 0.28 63.84 1.3725 ;
      RECT 63.775 0.8675 63.8625 1.0025 ;
      RECT 63.4 0.4875 63.465 1.14 ;
      RECT 63.4 0.6625 63.4825 0.7975 ;
      RECT 63.21 0.4875 63.275 1.14 ;
      RECT 63.1775 0.87 63.275 1.005 ;
      RECT 63.005 0.4875 63.07 1.14 ;
      RECT 63.005 0.87 63.1025 1.005 ;
      RECT 62.6425 1.25 62.7075 1.385 ;
      RECT 62.62 0.28 62.685 1.3725 ;
      RECT 62.055 0.265 62.12 1.3725 ;
      RECT 62.0325 0.725 62.12 0.86 ;
      RECT 61.6475 1.2375 61.735 1.3725 ;
      RECT 61.67 0.28 61.735 1.3725 ;
      RECT 61.465 0.4875 61.53 1.14 ;
      RECT 61.465 0.6825 61.5625 0.8175 ;
      RECT 61.275 0.4875 61.34 1.14 ;
      RECT 61.2575 0.8675 61.34 1.0025 ;
      RECT 61.09 0.4875 61.155 1.14 ;
      RECT 61.09 0.8675 61.1725 1.0025 ;
      RECT 60.9 0.485 60.965 1.14 ;
      RECT 60.8675 0.4675 60.9325 0.6025 ;
      RECT 60.515 0.28 60.58 1.3725 ;
      RECT 60.4925 0.6625 60.58 0.7975 ;
      RECT 60.31 0.28 60.375 1.3725 ;
      RECT 60.31 0.8675 60.3975 1.0025 ;
      RECT 59.935 0.4875 60 1.14 ;
      RECT 59.935 0.6625 60.0175 0.7975 ;
      RECT 59.745 0.4875 59.81 1.14 ;
      RECT 59.7125 0.87 59.81 1.005 ;
      RECT 59.54 0.4875 59.605 1.14 ;
      RECT 59.54 0.87 59.6375 1.005 ;
      RECT 59.1775 1.25 59.2425 1.385 ;
      RECT 59.155 0.28 59.22 1.3725 ;
      RECT 58.59 0.265 58.655 1.3725 ;
      RECT 58.5675 0.725 58.655 0.86 ;
      RECT 58.1825 1.2375 58.27 1.3725 ;
      RECT 58.205 0.28 58.27 1.3725 ;
      RECT 58 0.4875 58.065 1.14 ;
      RECT 58 0.6825 58.0975 0.8175 ;
      RECT 57.81 0.4875 57.875 1.14 ;
      RECT 57.7925 0.8675 57.875 1.0025 ;
      RECT 57.625 0.4875 57.69 1.14 ;
      RECT 57.625 0.8675 57.7075 1.0025 ;
      RECT 57.435 0.485 57.5 1.14 ;
      RECT 57.4025 0.4675 57.4675 0.6025 ;
      RECT 57.05 0.28 57.115 1.3725 ;
      RECT 57.0275 0.6625 57.115 0.7975 ;
      RECT 56.845 0.28 56.91 1.3725 ;
      RECT 56.845 0.8675 56.9325 1.0025 ;
      RECT 56.47 0.4875 56.535 1.14 ;
      RECT 56.47 0.6625 56.5525 0.7975 ;
      RECT 56.28 0.4875 56.345 1.14 ;
      RECT 56.2475 0.87 56.345 1.005 ;
      RECT 56.075 0.4875 56.14 1.14 ;
      RECT 56.075 0.87 56.1725 1.005 ;
      RECT 55.7125 1.25 55.7775 1.385 ;
      RECT 55.69 0.28 55.755 1.3725 ;
      RECT 55.125 0.265 55.19 1.3725 ;
      RECT 55.1025 0.725 55.19 0.86 ;
      RECT 54.7175 1.2375 54.805 1.3725 ;
      RECT 54.74 0.28 54.805 1.3725 ;
      RECT 54.535 0.4875 54.6 1.14 ;
      RECT 54.535 0.6825 54.6325 0.8175 ;
      RECT 54.345 0.4875 54.41 1.14 ;
      RECT 54.3275 0.8675 54.41 1.0025 ;
      RECT 54.16 0.4875 54.225 1.14 ;
      RECT 54.16 0.8675 54.2425 1.0025 ;
      RECT 53.97 0.485 54.035 1.14 ;
      RECT 53.9375 0.4675 54.0025 0.6025 ;
      RECT 53.585 0.28 53.65 1.3725 ;
      RECT 53.5625 0.6625 53.65 0.7975 ;
      RECT 53.38 0.28 53.445 1.3725 ;
      RECT 53.38 0.8675 53.4675 1.0025 ;
      RECT 53.005 0.4875 53.07 1.14 ;
      RECT 53.005 0.6625 53.0875 0.7975 ;
      RECT 52.815 0.4875 52.88 1.14 ;
      RECT 52.7825 0.87 52.88 1.005 ;
      RECT 52.61 0.4875 52.675 1.14 ;
      RECT 52.61 0.87 52.7075 1.005 ;
      RECT 52.2475 1.25 52.3125 1.385 ;
      RECT 52.225 0.28 52.29 1.3725 ;
      RECT 51.66 0.265 51.725 1.3725 ;
      RECT 51.6375 0.725 51.725 0.86 ;
      RECT 51.2525 1.2375 51.34 1.3725 ;
      RECT 51.275 0.28 51.34 1.3725 ;
      RECT 51.07 0.4875 51.135 1.14 ;
      RECT 51.07 0.6825 51.1675 0.8175 ;
      RECT 50.88 0.4875 50.945 1.14 ;
      RECT 50.8625 0.8675 50.945 1.0025 ;
      RECT 50.695 0.4875 50.76 1.14 ;
      RECT 50.695 0.8675 50.7775 1.0025 ;
      RECT 50.505 0.485 50.57 1.14 ;
      RECT 50.4725 0.4675 50.5375 0.6025 ;
      RECT 50.12 0.28 50.185 1.3725 ;
      RECT 50.0975 0.6625 50.185 0.7975 ;
      RECT 49.915 0.28 49.98 1.3725 ;
      RECT 49.915 0.8675 50.0025 1.0025 ;
      RECT 49.54 0.4875 49.605 1.14 ;
      RECT 49.54 0.6625 49.6225 0.7975 ;
      RECT 49.35 0.4875 49.415 1.14 ;
      RECT 49.3175 0.87 49.415 1.005 ;
      RECT 49.145 0.4875 49.21 1.14 ;
      RECT 49.145 0.87 49.2425 1.005 ;
      RECT 48.7825 1.25 48.8475 1.385 ;
      RECT 48.76 0.28 48.825 1.3725 ;
      RECT 48.195 0.265 48.26 1.3725 ;
      RECT 48.1725 0.725 48.26 0.86 ;
      RECT 47.7875 1.2375 47.875 1.3725 ;
      RECT 47.81 0.28 47.875 1.3725 ;
      RECT 47.605 0.4875 47.67 1.14 ;
      RECT 47.605 0.6825 47.7025 0.8175 ;
      RECT 47.415 0.4875 47.48 1.14 ;
      RECT 47.3975 0.8675 47.48 1.0025 ;
      RECT 47.23 0.4875 47.295 1.14 ;
      RECT 47.23 0.8675 47.3125 1.0025 ;
      RECT 47.04 0.485 47.105 1.14 ;
      RECT 47.0075 0.4675 47.0725 0.6025 ;
      RECT 46.655 0.28 46.72 1.3725 ;
      RECT 46.6325 0.6625 46.72 0.7975 ;
      RECT 46.45 0.28 46.515 1.3725 ;
      RECT 46.45 0.8675 46.5375 1.0025 ;
      RECT 46.075 0.4875 46.14 1.14 ;
      RECT 46.075 0.6625 46.1575 0.7975 ;
      RECT 45.885 0.4875 45.95 1.14 ;
      RECT 45.8525 0.87 45.95 1.005 ;
      RECT 45.68 0.4875 45.745 1.14 ;
      RECT 45.68 0.87 45.7775 1.005 ;
      RECT 45.3175 1.25 45.3825 1.385 ;
      RECT 45.295 0.28 45.36 1.3725 ;
      RECT 44.73 0.265 44.795 1.3725 ;
      RECT 44.7075 0.725 44.795 0.86 ;
      RECT 44.3225 1.2375 44.41 1.3725 ;
      RECT 44.345 0.28 44.41 1.3725 ;
      RECT 44.14 0.4875 44.205 1.14 ;
      RECT 44.14 0.6825 44.2375 0.8175 ;
      RECT 43.95 0.4875 44.015 1.14 ;
      RECT 43.9325 0.8675 44.015 1.0025 ;
      RECT 43.765 0.4875 43.83 1.14 ;
      RECT 43.765 0.8675 43.8475 1.0025 ;
      RECT 43.575 0.485 43.64 1.14 ;
      RECT 43.5425 0.4675 43.6075 0.6025 ;
      RECT 43.19 0.28 43.255 1.3725 ;
      RECT 43.1675 0.6625 43.255 0.7975 ;
      RECT 42.985 0.28 43.05 1.3725 ;
      RECT 42.985 0.8675 43.0725 1.0025 ;
      RECT 42.61 0.4875 42.675 1.14 ;
      RECT 42.61 0.6625 42.6925 0.7975 ;
      RECT 42.42 0.4875 42.485 1.14 ;
      RECT 42.3875 0.87 42.485 1.005 ;
      RECT 42.215 0.4875 42.28 1.14 ;
      RECT 42.215 0.87 42.3125 1.005 ;
      RECT 41.8525 1.25 41.9175 1.385 ;
      RECT 41.83 0.28 41.895 1.3725 ;
      RECT 41.265 0.265 41.33 1.3725 ;
      RECT 41.2425 0.725 41.33 0.86 ;
      RECT 40.8575 1.2375 40.945 1.3725 ;
      RECT 40.88 0.28 40.945 1.3725 ;
      RECT 40.675 0.4875 40.74 1.14 ;
      RECT 40.675 0.6825 40.7725 0.8175 ;
      RECT 40.485 0.4875 40.55 1.14 ;
      RECT 40.4675 0.8675 40.55 1.0025 ;
      RECT 40.3 0.4875 40.365 1.14 ;
      RECT 40.3 0.8675 40.3825 1.0025 ;
      RECT 40.11 0.485 40.175 1.14 ;
      RECT 40.0775 0.4675 40.1425 0.6025 ;
      RECT 39.725 0.28 39.79 1.3725 ;
      RECT 39.7025 0.6625 39.79 0.7975 ;
      RECT 39.52 0.28 39.585 1.3725 ;
      RECT 39.52 0.8675 39.6075 1.0025 ;
      RECT 39.145 0.4875 39.21 1.14 ;
      RECT 39.145 0.6625 39.2275 0.7975 ;
      RECT 38.955 0.4875 39.02 1.14 ;
      RECT 38.9225 0.87 39.02 1.005 ;
      RECT 38.75 0.4875 38.815 1.14 ;
      RECT 38.75 0.87 38.8475 1.005 ;
      RECT 38.3875 1.25 38.4525 1.385 ;
      RECT 38.365 0.28 38.43 1.3725 ;
      RECT 37.8 0.265 37.865 1.3725 ;
      RECT 37.7775 0.725 37.865 0.86 ;
      RECT 37.3925 1.2375 37.48 1.3725 ;
      RECT 37.415 0.28 37.48 1.3725 ;
      RECT 37.21 0.4875 37.275 1.14 ;
      RECT 37.21 0.6825 37.3075 0.8175 ;
      RECT 37.02 0.4875 37.085 1.14 ;
      RECT 37.0025 0.8675 37.085 1.0025 ;
      RECT 36.835 0.4875 36.9 1.14 ;
      RECT 36.835 0.8675 36.9175 1.0025 ;
      RECT 36.645 0.485 36.71 1.14 ;
      RECT 36.6125 0.4675 36.6775 0.6025 ;
      RECT 36.26 0.28 36.325 1.3725 ;
      RECT 36.2375 0.6625 36.325 0.7975 ;
      RECT 36.055 0.28 36.12 1.3725 ;
      RECT 36.055 0.8675 36.1425 1.0025 ;
      RECT 35.68 0.4875 35.745 1.14 ;
      RECT 35.68 0.6625 35.7625 0.7975 ;
      RECT 35.49 0.4875 35.555 1.14 ;
      RECT 35.4575 0.87 35.555 1.005 ;
      RECT 35.285 0.4875 35.35 1.14 ;
      RECT 35.285 0.87 35.3825 1.005 ;
      RECT 34.9225 1.25 34.9875 1.385 ;
      RECT 34.9 0.28 34.965 1.3725 ;
      RECT 34.335 0.265 34.4 1.3725 ;
      RECT 34.3125 0.725 34.4 0.86 ;
      RECT 33.9275 1.2375 34.015 1.3725 ;
      RECT 33.95 0.28 34.015 1.3725 ;
      RECT 33.745 0.4875 33.81 1.14 ;
      RECT 33.745 0.6825 33.8425 0.8175 ;
      RECT 33.555 0.4875 33.62 1.14 ;
      RECT 33.5375 0.8675 33.62 1.0025 ;
      RECT 33.37 0.4875 33.435 1.14 ;
      RECT 33.37 0.8675 33.4525 1.0025 ;
      RECT 33.18 0.485 33.245 1.14 ;
      RECT 33.1475 0.4675 33.2125 0.6025 ;
      RECT 32.795 0.28 32.86 1.3725 ;
      RECT 32.7725 0.6625 32.86 0.7975 ;
      RECT 32.59 0.28 32.655 1.3725 ;
      RECT 32.59 0.8675 32.6775 1.0025 ;
      RECT 32.215 0.4875 32.28 1.14 ;
      RECT 32.215 0.6625 32.2975 0.7975 ;
      RECT 32.025 0.4875 32.09 1.14 ;
      RECT 31.9925 0.87 32.09 1.005 ;
      RECT 31.82 0.4875 31.885 1.14 ;
      RECT 31.82 0.87 31.9175 1.005 ;
      RECT 31.4575 1.25 31.5225 1.385 ;
      RECT 31.435 0.28 31.5 1.3725 ;
      RECT 30.87 0.265 30.935 1.3725 ;
      RECT 30.8475 0.725 30.935 0.86 ;
      RECT 30.4625 1.2375 30.55 1.3725 ;
      RECT 30.485 0.28 30.55 1.3725 ;
      RECT 30.28 0.4875 30.345 1.14 ;
      RECT 30.28 0.6825 30.3775 0.8175 ;
      RECT 30.09 0.4875 30.155 1.14 ;
      RECT 30.0725 0.8675 30.155 1.0025 ;
      RECT 29.905 0.4875 29.97 1.14 ;
      RECT 29.905 0.8675 29.9875 1.0025 ;
      RECT 29.715 0.485 29.78 1.14 ;
      RECT 29.6825 0.4675 29.7475 0.6025 ;
      RECT 29.33 0.28 29.395 1.3725 ;
      RECT 29.3075 0.6625 29.395 0.7975 ;
      RECT 29.125 0.28 29.19 1.3725 ;
      RECT 29.125 0.8675 29.2125 1.0025 ;
      RECT 28.75 0.4875 28.815 1.14 ;
      RECT 28.75 0.6625 28.8325 0.7975 ;
      RECT 28.56 0.4875 28.625 1.14 ;
      RECT 28.5275 0.87 28.625 1.005 ;
      RECT 28.355 0.4875 28.42 1.14 ;
      RECT 28.355 0.87 28.4525 1.005 ;
      RECT 27.9925 1.25 28.0575 1.385 ;
      RECT 27.97 0.28 28.035 1.3725 ;
      RECT 27.405 0.265 27.47 1.3725 ;
      RECT 27.3825 0.725 27.47 0.86 ;
      RECT 26.9975 1.2375 27.085 1.3725 ;
      RECT 27.02 0.28 27.085 1.3725 ;
      RECT 26.815 0.4875 26.88 1.14 ;
      RECT 26.815 0.6825 26.9125 0.8175 ;
      RECT 26.625 0.4875 26.69 1.14 ;
      RECT 26.6075 0.8675 26.69 1.0025 ;
      RECT 26.44 0.4875 26.505 1.14 ;
      RECT 26.44 0.8675 26.5225 1.0025 ;
      RECT 26.25 0.485 26.315 1.14 ;
      RECT 26.2175 0.4675 26.2825 0.6025 ;
      RECT 25.865 0.28 25.93 1.3725 ;
      RECT 25.8425 0.6625 25.93 0.7975 ;
      RECT 25.66 0.28 25.725 1.3725 ;
      RECT 25.66 0.8675 25.7475 1.0025 ;
      RECT 25.285 0.4875 25.35 1.14 ;
      RECT 25.285 0.6625 25.3675 0.7975 ;
      RECT 25.095 0.4875 25.16 1.14 ;
      RECT 25.0625 0.87 25.16 1.005 ;
      RECT 24.89 0.4875 24.955 1.14 ;
      RECT 24.89 0.87 24.9875 1.005 ;
      RECT 24.5275 1.25 24.5925 1.385 ;
      RECT 24.505 0.28 24.57 1.3725 ;
      RECT 23.94 0.265 24.005 1.3725 ;
      RECT 23.9175 0.725 24.005 0.86 ;
      RECT 23.5325 1.2375 23.62 1.3725 ;
      RECT 23.555 0.28 23.62 1.3725 ;
      RECT 23.35 0.4875 23.415 1.14 ;
      RECT 23.35 0.6825 23.4475 0.8175 ;
      RECT 23.16 0.4875 23.225 1.14 ;
      RECT 23.1425 0.8675 23.225 1.0025 ;
      RECT 22.975 0.4875 23.04 1.14 ;
      RECT 22.975 0.8675 23.0575 1.0025 ;
      RECT 22.785 0.485 22.85 1.14 ;
      RECT 22.7525 0.4675 22.8175 0.6025 ;
      RECT 22.4 0.28 22.465 1.3725 ;
      RECT 22.3775 0.6625 22.465 0.7975 ;
      RECT 22.195 0.28 22.26 1.3725 ;
      RECT 22.195 0.8675 22.2825 1.0025 ;
      RECT 21.82 0.4875 21.885 1.14 ;
      RECT 21.82 0.6625 21.9025 0.7975 ;
      RECT 21.63 0.4875 21.695 1.14 ;
      RECT 21.5975 0.87 21.695 1.005 ;
      RECT 21.425 0.4875 21.49 1.14 ;
      RECT 21.425 0.87 21.5225 1.005 ;
      RECT 21.0625 1.25 21.1275 1.385 ;
      RECT 21.04 0.28 21.105 1.3725 ;
      RECT 20.475 0.265 20.54 1.3725 ;
      RECT 20.4525 0.725 20.54 0.86 ;
      RECT 20.0675 1.2375 20.155 1.3725 ;
      RECT 20.09 0.28 20.155 1.3725 ;
      RECT 19.885 0.4875 19.95 1.14 ;
      RECT 19.885 0.6825 19.9825 0.8175 ;
      RECT 19.695 0.4875 19.76 1.14 ;
      RECT 19.6775 0.8675 19.76 1.0025 ;
      RECT 19.51 0.4875 19.575 1.14 ;
      RECT 19.51 0.8675 19.5925 1.0025 ;
      RECT 19.32 0.485 19.385 1.14 ;
      RECT 19.2875 0.4675 19.3525 0.6025 ;
      RECT 18.935 0.28 19 1.3725 ;
      RECT 18.9125 0.6625 19 0.7975 ;
      RECT 18.73 0.28 18.795 1.3725 ;
      RECT 18.73 0.8675 18.8175 1.0025 ;
      RECT 18.355 0.4875 18.42 1.14 ;
      RECT 18.355 0.6625 18.4375 0.7975 ;
      RECT 18.165 0.4875 18.23 1.14 ;
      RECT 18.1325 0.87 18.23 1.005 ;
      RECT 17.96 0.4875 18.025 1.14 ;
      RECT 17.96 0.87 18.0575 1.005 ;
      RECT 17.5975 1.25 17.6625 1.385 ;
      RECT 17.575 0.28 17.64 1.3725 ;
      RECT 17.01 0.265 17.075 1.3725 ;
      RECT 16.9875 0.725 17.075 0.86 ;
      RECT 16.6025 1.2375 16.69 1.3725 ;
      RECT 16.625 0.28 16.69 1.3725 ;
      RECT 16.42 0.4875 16.485 1.14 ;
      RECT 16.42 0.6825 16.5175 0.8175 ;
      RECT 16.23 0.4875 16.295 1.14 ;
      RECT 16.2125 0.8675 16.295 1.0025 ;
      RECT 16.045 0.4875 16.11 1.14 ;
      RECT 16.045 0.8675 16.1275 1.0025 ;
      RECT 15.855 0.485 15.92 1.14 ;
      RECT 15.8225 0.4675 15.8875 0.6025 ;
      RECT 15.47 0.28 15.535 1.3725 ;
      RECT 15.4475 0.6625 15.535 0.7975 ;
      RECT 15.265 0.28 15.33 1.3725 ;
      RECT 15.265 0.8675 15.3525 1.0025 ;
      RECT 14.89 0.4875 14.955 1.14 ;
      RECT 14.89 0.6625 14.9725 0.7975 ;
      RECT 14.7 0.4875 14.765 1.14 ;
      RECT 14.6675 0.87 14.765 1.005 ;
      RECT 14.495 0.4875 14.56 1.14 ;
      RECT 14.495 0.87 14.5925 1.005 ;
      RECT 14.1325 1.25 14.1975 1.385 ;
      RECT 14.11 0.28 14.175 1.3725 ;
      RECT 13.545 0.265 13.61 1.3725 ;
      RECT 13.5225 0.725 13.61 0.86 ;
      RECT 13.1375 1.2375 13.225 1.3725 ;
      RECT 13.16 0.28 13.225 1.3725 ;
      RECT 12.955 0.4875 13.02 1.14 ;
      RECT 12.955 0.6825 13.0525 0.8175 ;
      RECT 12.765 0.4875 12.83 1.14 ;
      RECT 12.7475 0.8675 12.83 1.0025 ;
      RECT 12.58 0.4875 12.645 1.14 ;
      RECT 12.58 0.8675 12.6625 1.0025 ;
      RECT 12.39 0.485 12.455 1.14 ;
      RECT 12.3575 0.4675 12.4225 0.6025 ;
      RECT 12.005 0.28 12.07 1.3725 ;
      RECT 11.9825 0.6625 12.07 0.7975 ;
      RECT 11.8 0.28 11.865 1.3725 ;
      RECT 11.8 0.8675 11.8875 1.0025 ;
      RECT 11.425 0.4875 11.49 1.14 ;
      RECT 11.425 0.6625 11.5075 0.7975 ;
      RECT 11.235 0.4875 11.3 1.14 ;
      RECT 11.2025 0.87 11.3 1.005 ;
      RECT 11.03 0.4875 11.095 1.14 ;
      RECT 11.03 0.87 11.1275 1.005 ;
      RECT 10.6675 1.25 10.7325 1.385 ;
      RECT 10.645 0.28 10.71 1.3725 ;
      RECT 10.08 0.265 10.145 1.3725 ;
      RECT 10.0575 0.725 10.145 0.86 ;
      RECT 9.6725 1.2375 9.76 1.3725 ;
      RECT 9.695 0.28 9.76 1.3725 ;
      RECT 9.49 0.4875 9.555 1.14 ;
      RECT 9.49 0.6825 9.5875 0.8175 ;
      RECT 9.3 0.4875 9.365 1.14 ;
      RECT 9.2825 0.8675 9.365 1.0025 ;
      RECT 9.115 0.4875 9.18 1.14 ;
      RECT 9.115 0.8675 9.1975 1.0025 ;
      RECT 8.925 0.485 8.99 1.14 ;
      RECT 8.8925 0.4675 8.9575 0.6025 ;
      RECT 8.54 0.28 8.605 1.3725 ;
      RECT 8.5175 0.6625 8.605 0.7975 ;
      RECT 8.335 0.28 8.4 1.3725 ;
      RECT 8.335 0.8675 8.4225 1.0025 ;
      RECT 7.96 0.4875 8.025 1.14 ;
      RECT 7.96 0.6625 8.0425 0.7975 ;
      RECT 7.77 0.4875 7.835 1.14 ;
      RECT 7.7375 0.87 7.835 1.005 ;
      RECT 7.565 0.4875 7.63 1.14 ;
      RECT 7.565 0.87 7.6625 1.005 ;
      RECT 7.2025 1.25 7.2675 1.385 ;
      RECT 7.18 0.28 7.245 1.3725 ;
      RECT 6.615 0.265 6.68 1.3725 ;
      RECT 6.5925 0.725 6.68 0.86 ;
      RECT 6.2075 1.2375 6.295 1.3725 ;
      RECT 6.23 0.28 6.295 1.3725 ;
      RECT 6.025 0.4875 6.09 1.14 ;
      RECT 6.025 0.6825 6.1225 0.8175 ;
      RECT 5.835 0.4875 5.9 1.14 ;
      RECT 5.8175 0.8675 5.9 1.0025 ;
      RECT 5.65 0.4875 5.715 1.14 ;
      RECT 5.65 0.8675 5.7325 1.0025 ;
      RECT 5.46 0.485 5.525 1.14 ;
      RECT 5.4275 0.4675 5.4925 0.6025 ;
      RECT 5.075 0.28 5.14 1.3725 ;
      RECT 5.0525 0.6625 5.14 0.7975 ;
      RECT 4.87 0.28 4.935 1.3725 ;
      RECT 4.87 0.8675 4.9575 1.0025 ;
      RECT 4.495 0.4875 4.56 1.14 ;
      RECT 4.495 0.6625 4.5775 0.7975 ;
      RECT 4.305 0.4875 4.37 1.14 ;
      RECT 4.2725 0.87 4.37 1.005 ;
      RECT 4.1 0.4875 4.165 1.14 ;
      RECT 4.1 0.87 4.1975 1.005 ;
      RECT 3.7375 1.25 3.8025 1.385 ;
      RECT 3.715 0.28 3.78 1.3725 ;
      RECT 3.15 0.265 3.215 1.3725 ;
      RECT 3.1275 0.725 3.215 0.86 ;
      RECT 2.7425 1.2375 2.83 1.3725 ;
      RECT 2.765 0.28 2.83 1.3725 ;
      RECT 2.56 0.4875 2.625 1.14 ;
      RECT 2.56 0.6825 2.6575 0.8175 ;
      RECT 2.37 0.4875 2.435 1.14 ;
      RECT 2.3525 0.8675 2.435 1.0025 ;
      RECT 2.185 0.4875 2.25 1.14 ;
      RECT 2.185 0.8675 2.2675 1.0025 ;
      RECT 1.995 0.485 2.06 1.14 ;
      RECT 1.9625 0.4675 2.0275 0.6025 ;
      RECT 1.61 0.28 1.675 1.3725 ;
      RECT 1.5875 0.6625 1.675 0.7975 ;
      RECT 1.405 0.28 1.47 1.3725 ;
      RECT 1.405 0.8675 1.4925 1.0025 ;
      RECT 1.03 0.4875 1.095 1.14 ;
      RECT 1.03 0.6625 1.1125 0.7975 ;
      RECT 0.84 0.4875 0.905 1.14 ;
      RECT 0.8075 0.87 0.905 1.005 ;
      RECT 0.635 0.4875 0.7 1.14 ;
      RECT 0.635 0.87 0.7325 1.005 ;
      RECT 0.2725 1.25 0.3375 1.385 ;
      RECT 0.25 0.28 0.315 1.3725 ;
      RECT 115.17 1.03 115.235 1.165 ;
      RECT 114.845 0.265 114.91 1.355 ;
      RECT 114.715 0.405 114.78 0.54 ;
      RECT 114.715 0.96 114.78 1.095 ;
      RECT 114.585 0.265 114.65 1.355 ;
      RECT 114.455 0.405 114.52 0.54 ;
      RECT 114.455 1.015 114.52 1.15 ;
      RECT 114.1325 0.7075 114.2025 0.8425 ;
      RECT 113.98 0.265 114.045 1.3425 ;
      RECT 113.7375 0.47 113.8025 0.605 ;
      RECT 113.2825 0.47 113.3475 0.605 ;
      RECT 113.04 0.265 113.105 1.3425 ;
      RECT 112.8825 0.4525 112.9525 0.5875 ;
      RECT 112.565 0.405 112.63 0.54 ;
      RECT 112.565 1.015 112.63 1.15 ;
      RECT 112.435 0.265 112.5 1.355 ;
      RECT 112.305 0.405 112.37 0.54 ;
      RECT 112.305 0.96 112.37 1.095 ;
      RECT 112.175 0.265 112.24 1.355 ;
      RECT 111.85 1.03 111.915 1.165 ;
      RECT 111.3575 0.455 111.4225 0.59 ;
      RECT 110.9725 0.68 111.0375 0.815 ;
      RECT 109.8425 1.27 109.9775 1.335 ;
      RECT 109.4725 1.315 109.6075 1.38 ;
      RECT 109.1825 0.8675 109.2475 1.0025 ;
      RECT 108.6625 0.8675 108.7275 1.0025 ;
      RECT 108.3475 0.2825 108.4125 0.4175 ;
      RECT 107.9175 1.2725 108.0525 1.3375 ;
      RECT 106.3775 1.27 106.5125 1.335 ;
      RECT 106.0075 1.315 106.1425 1.38 ;
      RECT 105.7175 0.8675 105.7825 1.0025 ;
      RECT 105.1975 0.8675 105.2625 1.0025 ;
      RECT 104.8825 0.2825 104.9475 0.4175 ;
      RECT 104.4525 1.2725 104.5875 1.3375 ;
      RECT 102.9125 1.27 103.0475 1.335 ;
      RECT 102.5425 1.315 102.6775 1.38 ;
      RECT 102.2525 0.8675 102.3175 1.0025 ;
      RECT 101.7325 0.8675 101.7975 1.0025 ;
      RECT 101.4175 0.2825 101.4825 0.4175 ;
      RECT 100.9875 1.2725 101.1225 1.3375 ;
      RECT 99.4475 1.27 99.5825 1.335 ;
      RECT 99.0775 1.315 99.2125 1.38 ;
      RECT 98.7875 0.8675 98.8525 1.0025 ;
      RECT 98.2675 0.8675 98.3325 1.0025 ;
      RECT 97.9525 0.2825 98.0175 0.4175 ;
      RECT 97.5225 1.2725 97.6575 1.3375 ;
      RECT 95.9825 1.27 96.1175 1.335 ;
      RECT 95.6125 1.315 95.7475 1.38 ;
      RECT 95.3225 0.8675 95.3875 1.0025 ;
      RECT 94.8025 0.8675 94.8675 1.0025 ;
      RECT 94.4875 0.2825 94.5525 0.4175 ;
      RECT 94.0575 1.2725 94.1925 1.3375 ;
      RECT 92.5175 1.27 92.6525 1.335 ;
      RECT 92.1475 1.315 92.2825 1.38 ;
      RECT 91.8575 0.8675 91.9225 1.0025 ;
      RECT 91.3375 0.8675 91.4025 1.0025 ;
      RECT 91.0225 0.2825 91.0875 0.4175 ;
      RECT 90.5925 1.2725 90.7275 1.3375 ;
      RECT 89.0525 1.27 89.1875 1.335 ;
      RECT 88.6825 1.315 88.8175 1.38 ;
      RECT 88.3925 0.8675 88.4575 1.0025 ;
      RECT 87.8725 0.8675 87.9375 1.0025 ;
      RECT 87.5575 0.2825 87.6225 0.4175 ;
      RECT 87.1275 1.2725 87.2625 1.3375 ;
      RECT 85.5875 1.27 85.7225 1.335 ;
      RECT 85.2175 1.315 85.3525 1.38 ;
      RECT 84.9275 0.8675 84.9925 1.0025 ;
      RECT 84.4075 0.8675 84.4725 1.0025 ;
      RECT 84.0925 0.2825 84.1575 0.4175 ;
      RECT 83.6625 1.2725 83.7975 1.3375 ;
      RECT 82.1225 1.27 82.2575 1.335 ;
      RECT 81.7525 1.315 81.8875 1.38 ;
      RECT 81.4625 0.8675 81.5275 1.0025 ;
      RECT 80.9425 0.8675 81.0075 1.0025 ;
      RECT 80.6275 0.2825 80.6925 0.4175 ;
      RECT 80.1975 1.2725 80.3325 1.3375 ;
      RECT 78.6575 1.27 78.7925 1.335 ;
      RECT 78.2875 1.315 78.4225 1.38 ;
      RECT 77.9975 0.8675 78.0625 1.0025 ;
      RECT 77.4775 0.8675 77.5425 1.0025 ;
      RECT 77.1625 0.2825 77.2275 0.4175 ;
      RECT 76.7325 1.2725 76.8675 1.3375 ;
      RECT 75.1925 1.27 75.3275 1.335 ;
      RECT 74.8225 1.315 74.9575 1.38 ;
      RECT 74.5325 0.8675 74.5975 1.0025 ;
      RECT 74.0125 0.8675 74.0775 1.0025 ;
      RECT 73.6975 0.2825 73.7625 0.4175 ;
      RECT 73.2675 1.2725 73.4025 1.3375 ;
      RECT 71.7275 1.27 71.8625 1.335 ;
      RECT 71.3575 1.315 71.4925 1.38 ;
      RECT 71.0675 0.8675 71.1325 1.0025 ;
      RECT 70.5475 0.8675 70.6125 1.0025 ;
      RECT 70.2325 0.2825 70.2975 0.4175 ;
      RECT 69.8025 1.2725 69.9375 1.3375 ;
      RECT 68.2625 1.27 68.3975 1.335 ;
      RECT 67.8925 1.315 68.0275 1.38 ;
      RECT 67.6025 0.8675 67.6675 1.0025 ;
      RECT 67.0825 0.8675 67.1475 1.0025 ;
      RECT 66.7675 0.2825 66.8325 0.4175 ;
      RECT 66.3375 1.2725 66.4725 1.3375 ;
      RECT 64.7975 1.27 64.9325 1.335 ;
      RECT 64.4275 1.315 64.5625 1.38 ;
      RECT 64.1375 0.8675 64.2025 1.0025 ;
      RECT 63.6175 0.8675 63.6825 1.0025 ;
      RECT 63.3025 0.2825 63.3675 0.4175 ;
      RECT 62.8725 1.2725 63.0075 1.3375 ;
      RECT 61.3325 1.27 61.4675 1.335 ;
      RECT 60.9625 1.315 61.0975 1.38 ;
      RECT 60.6725 0.8675 60.7375 1.0025 ;
      RECT 60.1525 0.8675 60.2175 1.0025 ;
      RECT 59.8375 0.2825 59.9025 0.4175 ;
      RECT 59.4075 1.2725 59.5425 1.3375 ;
      RECT 57.8675 1.27 58.0025 1.335 ;
      RECT 57.4975 1.315 57.6325 1.38 ;
      RECT 57.2075 0.8675 57.2725 1.0025 ;
      RECT 56.6875 0.8675 56.7525 1.0025 ;
      RECT 56.3725 0.2825 56.4375 0.4175 ;
      RECT 55.9425 1.2725 56.0775 1.3375 ;
      RECT 54.4025 1.27 54.5375 1.335 ;
      RECT 54.0325 1.315 54.1675 1.38 ;
      RECT 53.7425 0.8675 53.8075 1.0025 ;
      RECT 53.2225 0.8675 53.2875 1.0025 ;
      RECT 52.9075 0.2825 52.9725 0.4175 ;
      RECT 52.4775 1.2725 52.6125 1.3375 ;
      RECT 50.9375 1.27 51.0725 1.335 ;
      RECT 50.5675 1.315 50.7025 1.38 ;
      RECT 50.2775 0.8675 50.3425 1.0025 ;
      RECT 49.7575 0.8675 49.8225 1.0025 ;
      RECT 49.4425 0.2825 49.5075 0.4175 ;
      RECT 49.0125 1.2725 49.1475 1.3375 ;
      RECT 47.4725 1.27 47.6075 1.335 ;
      RECT 47.1025 1.315 47.2375 1.38 ;
      RECT 46.8125 0.8675 46.8775 1.0025 ;
      RECT 46.2925 0.8675 46.3575 1.0025 ;
      RECT 45.9775 0.2825 46.0425 0.4175 ;
      RECT 45.5475 1.2725 45.6825 1.3375 ;
      RECT 44.0075 1.27 44.1425 1.335 ;
      RECT 43.6375 1.315 43.7725 1.38 ;
      RECT 43.3475 0.8675 43.4125 1.0025 ;
      RECT 42.8275 0.8675 42.8925 1.0025 ;
      RECT 42.5125 0.2825 42.5775 0.4175 ;
      RECT 42.0825 1.2725 42.2175 1.3375 ;
      RECT 40.5425 1.27 40.6775 1.335 ;
      RECT 40.1725 1.315 40.3075 1.38 ;
      RECT 39.8825 0.8675 39.9475 1.0025 ;
      RECT 39.3625 0.8675 39.4275 1.0025 ;
      RECT 39.0475 0.2825 39.1125 0.4175 ;
      RECT 38.6175 1.2725 38.7525 1.3375 ;
      RECT 37.0775 1.27 37.2125 1.335 ;
      RECT 36.7075 1.315 36.8425 1.38 ;
      RECT 36.4175 0.8675 36.4825 1.0025 ;
      RECT 35.8975 0.8675 35.9625 1.0025 ;
      RECT 35.5825 0.2825 35.6475 0.4175 ;
      RECT 35.1525 1.2725 35.2875 1.3375 ;
      RECT 33.6125 1.27 33.7475 1.335 ;
      RECT 33.2425 1.315 33.3775 1.38 ;
      RECT 32.9525 0.8675 33.0175 1.0025 ;
      RECT 32.4325 0.8675 32.4975 1.0025 ;
      RECT 32.1175 0.2825 32.1825 0.4175 ;
      RECT 31.6875 1.2725 31.8225 1.3375 ;
      RECT 30.1475 1.27 30.2825 1.335 ;
      RECT 29.7775 1.315 29.9125 1.38 ;
      RECT 29.4875 0.8675 29.5525 1.0025 ;
      RECT 28.9675 0.8675 29.0325 1.0025 ;
      RECT 28.6525 0.2825 28.7175 0.4175 ;
      RECT 28.2225 1.2725 28.3575 1.3375 ;
      RECT 26.6825 1.27 26.8175 1.335 ;
      RECT 26.3125 1.315 26.4475 1.38 ;
      RECT 26.0225 0.8675 26.0875 1.0025 ;
      RECT 25.5025 0.8675 25.5675 1.0025 ;
      RECT 25.1875 0.2825 25.2525 0.4175 ;
      RECT 24.7575 1.2725 24.8925 1.3375 ;
      RECT 23.2175 1.27 23.3525 1.335 ;
      RECT 22.8475 1.315 22.9825 1.38 ;
      RECT 22.5575 0.8675 22.6225 1.0025 ;
      RECT 22.0375 0.8675 22.1025 1.0025 ;
      RECT 21.7225 0.2825 21.7875 0.4175 ;
      RECT 21.2925 1.2725 21.4275 1.3375 ;
      RECT 19.7525 1.27 19.8875 1.335 ;
      RECT 19.3825 1.315 19.5175 1.38 ;
      RECT 19.0925 0.8675 19.1575 1.0025 ;
      RECT 18.5725 0.8675 18.6375 1.0025 ;
      RECT 18.2575 0.2825 18.3225 0.4175 ;
      RECT 17.8275 1.2725 17.9625 1.3375 ;
      RECT 16.2875 1.27 16.4225 1.335 ;
      RECT 15.9175 1.315 16.0525 1.38 ;
      RECT 15.6275 0.8675 15.6925 1.0025 ;
      RECT 15.1075 0.8675 15.1725 1.0025 ;
      RECT 14.7925 0.2825 14.8575 0.4175 ;
      RECT 14.3625 1.2725 14.4975 1.3375 ;
      RECT 12.8225 1.27 12.9575 1.335 ;
      RECT 12.4525 1.315 12.5875 1.38 ;
      RECT 12.1625 0.8675 12.2275 1.0025 ;
      RECT 11.6425 0.8675 11.7075 1.0025 ;
      RECT 11.3275 0.2825 11.3925 0.4175 ;
      RECT 10.8975 1.2725 11.0325 1.3375 ;
      RECT 9.3575 1.27 9.4925 1.335 ;
      RECT 8.9875 1.315 9.1225 1.38 ;
      RECT 8.6975 0.8675 8.7625 1.0025 ;
      RECT 8.1775 0.8675 8.2425 1.0025 ;
      RECT 7.8625 0.2825 7.9275 0.4175 ;
      RECT 7.4325 1.2725 7.5675 1.3375 ;
      RECT 5.8925 1.27 6.0275 1.335 ;
      RECT 5.5225 1.315 5.6575 1.38 ;
      RECT 5.2325 0.8675 5.2975 1.0025 ;
      RECT 4.7125 0.8675 4.7775 1.0025 ;
      RECT 4.3975 0.2825 4.4625 0.4175 ;
      RECT 3.9675 1.2725 4.1025 1.3375 ;
      RECT 2.4275 1.27 2.5625 1.335 ;
      RECT 2.0575 1.315 2.1925 1.38 ;
      RECT 1.7675 0.8675 1.8325 1.0025 ;
      RECT 1.2475 0.8675 1.3125 1.0025 ;
      RECT 0.9325 0.2825 0.9975 0.4175 ;
      RECT 0.5025 1.2725 0.6375 1.3375 ;
    LAYER metal2 ;
      RECT 114.5825 1.3125 115.2325 1.3825 ;
      RECT 115.1625 1.03 115.2325 1.3825 ;
      RECT 114.5825 1.22 114.6525 1.3825 ;
      RECT 115.1625 1.03 115.2375 1.165 ;
      RECT 114.7125 0.96 114.7825 1.095 ;
      RECT 114.715 0.75 114.785 1.02 ;
      RECT 114.715 0.75 115.0425 0.82 ;
      RECT 114.9725 0.125 115.0425 0.82 ;
      RECT 114.425 0.405 114.5225 0.54 ;
      RECT 114.425 0.125 114.495 0.54 ;
      RECT 113.6 0.125 113.67 0.4 ;
      RECT 113.6 0.125 115.0425 0.195 ;
      RECT 113.9775 1.0375 114.0475 1.3425 ;
      RECT 114.4525 0.61 114.5225 1.15 ;
      RECT 113.9775 1.0375 114.5225 1.1075 ;
      RECT 114.4525 0.61 114.78 0.68 ;
      RECT 114.71 0.4275 114.78 0.68 ;
      RECT 114.7125 0.405 114.7825 0.54 ;
      RECT 113.9775 0.4725 114.0475 0.6075 ;
      RECT 113.735 0.47 113.805 0.605 ;
      RECT 113.73 0.5 114.05 0.57 ;
      RECT 112.3025 0.96 112.3725 1.095 ;
      RECT 112.3 0.75 112.37 1.02 ;
      RECT 112.0425 0.75 112.37 0.82 ;
      RECT 112.0425 0.125 112.1125 0.82 ;
      RECT 112.5625 0.405 112.66 0.54 ;
      RECT 112.59 0.125 112.66 0.54 ;
      RECT 113.415 0.125 113.485 0.4 ;
      RECT 112.0425 0.125 113.485 0.195 ;
      RECT 113.0375 0.4725 113.1075 0.6075 ;
      RECT 113.28 0.47 113.35 0.605 ;
      RECT 113.035 0.5 113.355 0.57 ;
      RECT 113.0375 1.0375 113.1075 1.3425 ;
      RECT 112.5625 0.61 112.6325 1.15 ;
      RECT 112.5625 1.0375 113.1075 1.1075 ;
      RECT 112.305 0.61 112.6325 0.68 ;
      RECT 112.305 0.4275 112.375 0.68 ;
      RECT 112.3025 0.405 112.3725 0.54 ;
      RECT 111.8525 1.32 112.5025 1.39 ;
      RECT 112.4325 1.22 112.5025 1.39 ;
      RECT 111.8525 1.03 111.9225 1.39 ;
      RECT 111.8475 1.03 111.9225 1.165 ;
      RECT 109.5025 1.455 110.63 1.525 ;
      RECT 110.56 0.725 110.63 1.525 ;
      RECT 109.5025 1.3125 109.5725 1.525 ;
      RECT 109.4725 1.3125 109.6075 1.3825 ;
      RECT 110.54 0.725 110.63 0.86 ;
      RECT 110.155 1.2375 110.225 1.3725 ;
      RECT 109.8425 1.2675 110.225 1.3375 ;
      RECT 109.765 0.8675 109.835 1.0025 ;
      RECT 109.615 0.8675 109.685 1.0025 ;
      RECT 109.18 0.8675 109.25 1.0025 ;
      RECT 108.84 0.8675 108.91 1.0025 ;
      RECT 108.84 0.9025 109.835 0.9725 ;
      RECT 109 0.6625 109.07 0.7975 ;
      RECT 108.46 0.6625 108.53 0.7975 ;
      RECT 108.46 0.695 109.07 0.765 ;
      RECT 108.22 0.87 108.29 1.005 ;
      RECT 108.08 0.87 108.15 1.005 ;
      RECT 108.66 0.8675 108.73 1.0025 ;
      RECT 108.08 0.9025 108.7325 0.9725 ;
      RECT 107.685 1.225 107.755 1.385 ;
      RECT 107.9175 1.225 108.0525 1.34 ;
      RECT 107.6875 0.5425 107.7575 1.32 ;
      RECT 107.685 1.225 108.0525 1.295 ;
      RECT 107.6875 0.5425 108.2 0.6125 ;
      RECT 108.13 0.3375 108.2 0.6125 ;
      RECT 108.345 0.2825 108.415 0.4175 ;
      RECT 108.13 0.3375 108.4175 0.4075 ;
      RECT 106.0375 1.455 107.165 1.525 ;
      RECT 107.095 0.725 107.165 1.525 ;
      RECT 106.0375 1.3125 106.1075 1.525 ;
      RECT 106.0075 1.3125 106.1425 1.3825 ;
      RECT 107.075 0.725 107.165 0.86 ;
      RECT 106.69 1.2375 106.76 1.3725 ;
      RECT 106.3775 1.2675 106.76 1.3375 ;
      RECT 106.3 0.8675 106.37 1.0025 ;
      RECT 106.15 0.8675 106.22 1.0025 ;
      RECT 105.715 0.8675 105.785 1.0025 ;
      RECT 105.375 0.8675 105.445 1.0025 ;
      RECT 105.375 0.9025 106.37 0.9725 ;
      RECT 105.535 0.6625 105.605 0.7975 ;
      RECT 104.995 0.6625 105.065 0.7975 ;
      RECT 104.995 0.695 105.605 0.765 ;
      RECT 104.755 0.87 104.825 1.005 ;
      RECT 104.615 0.87 104.685 1.005 ;
      RECT 105.195 0.8675 105.265 1.0025 ;
      RECT 104.615 0.9025 105.2675 0.9725 ;
      RECT 104.22 1.225 104.29 1.385 ;
      RECT 104.4525 1.225 104.5875 1.34 ;
      RECT 104.2225 0.5425 104.2925 1.32 ;
      RECT 104.22 1.225 104.5875 1.295 ;
      RECT 104.2225 0.5425 104.735 0.6125 ;
      RECT 104.665 0.3375 104.735 0.6125 ;
      RECT 104.88 0.2825 104.95 0.4175 ;
      RECT 104.665 0.3375 104.9525 0.4075 ;
      RECT 102.5725 1.455 103.7 1.525 ;
      RECT 103.63 0.725 103.7 1.525 ;
      RECT 102.5725 1.3125 102.6425 1.525 ;
      RECT 102.5425 1.3125 102.6775 1.3825 ;
      RECT 103.61 0.725 103.7 0.86 ;
      RECT 103.225 1.2375 103.295 1.3725 ;
      RECT 102.9125 1.2675 103.295 1.3375 ;
      RECT 102.835 0.8675 102.905 1.0025 ;
      RECT 102.685 0.8675 102.755 1.0025 ;
      RECT 102.25 0.8675 102.32 1.0025 ;
      RECT 101.91 0.8675 101.98 1.0025 ;
      RECT 101.91 0.9025 102.905 0.9725 ;
      RECT 102.07 0.6625 102.14 0.7975 ;
      RECT 101.53 0.6625 101.6 0.7975 ;
      RECT 101.53 0.695 102.14 0.765 ;
      RECT 101.29 0.87 101.36 1.005 ;
      RECT 101.15 0.87 101.22 1.005 ;
      RECT 101.73 0.8675 101.8 1.0025 ;
      RECT 101.15 0.9025 101.8025 0.9725 ;
      RECT 100.755 1.225 100.825 1.385 ;
      RECT 100.9875 1.225 101.1225 1.34 ;
      RECT 100.7575 0.5425 100.8275 1.32 ;
      RECT 100.755 1.225 101.1225 1.295 ;
      RECT 100.7575 0.5425 101.27 0.6125 ;
      RECT 101.2 0.3375 101.27 0.6125 ;
      RECT 101.415 0.2825 101.485 0.4175 ;
      RECT 101.2 0.3375 101.4875 0.4075 ;
      RECT 99.1075 1.455 100.235 1.525 ;
      RECT 100.165 0.725 100.235 1.525 ;
      RECT 99.1075 1.3125 99.1775 1.525 ;
      RECT 99.0775 1.3125 99.2125 1.3825 ;
      RECT 100.145 0.725 100.235 0.86 ;
      RECT 99.76 1.2375 99.83 1.3725 ;
      RECT 99.4475 1.2675 99.83 1.3375 ;
      RECT 99.37 0.8675 99.44 1.0025 ;
      RECT 99.22 0.8675 99.29 1.0025 ;
      RECT 98.785 0.8675 98.855 1.0025 ;
      RECT 98.445 0.8675 98.515 1.0025 ;
      RECT 98.445 0.9025 99.44 0.9725 ;
      RECT 98.605 0.6625 98.675 0.7975 ;
      RECT 98.065 0.6625 98.135 0.7975 ;
      RECT 98.065 0.695 98.675 0.765 ;
      RECT 97.825 0.87 97.895 1.005 ;
      RECT 97.685 0.87 97.755 1.005 ;
      RECT 98.265 0.8675 98.335 1.0025 ;
      RECT 97.685 0.9025 98.3375 0.9725 ;
      RECT 97.29 1.225 97.36 1.385 ;
      RECT 97.5225 1.225 97.6575 1.34 ;
      RECT 97.2925 0.5425 97.3625 1.32 ;
      RECT 97.29 1.225 97.6575 1.295 ;
      RECT 97.2925 0.5425 97.805 0.6125 ;
      RECT 97.735 0.3375 97.805 0.6125 ;
      RECT 97.95 0.2825 98.02 0.4175 ;
      RECT 97.735 0.3375 98.0225 0.4075 ;
      RECT 95.6425 1.455 96.77 1.525 ;
      RECT 96.7 0.725 96.77 1.525 ;
      RECT 95.6425 1.3125 95.7125 1.525 ;
      RECT 95.6125 1.3125 95.7475 1.3825 ;
      RECT 96.68 0.725 96.77 0.86 ;
      RECT 96.295 1.2375 96.365 1.3725 ;
      RECT 95.9825 1.2675 96.365 1.3375 ;
      RECT 95.905 0.8675 95.975 1.0025 ;
      RECT 95.755 0.8675 95.825 1.0025 ;
      RECT 95.32 0.8675 95.39 1.0025 ;
      RECT 94.98 0.8675 95.05 1.0025 ;
      RECT 94.98 0.9025 95.975 0.9725 ;
      RECT 95.14 0.6625 95.21 0.7975 ;
      RECT 94.6 0.6625 94.67 0.7975 ;
      RECT 94.6 0.695 95.21 0.765 ;
      RECT 94.36 0.87 94.43 1.005 ;
      RECT 94.22 0.87 94.29 1.005 ;
      RECT 94.8 0.8675 94.87 1.0025 ;
      RECT 94.22 0.9025 94.8725 0.9725 ;
      RECT 93.825 1.225 93.895 1.385 ;
      RECT 94.0575 1.225 94.1925 1.34 ;
      RECT 93.8275 0.5425 93.8975 1.32 ;
      RECT 93.825 1.225 94.1925 1.295 ;
      RECT 93.8275 0.5425 94.34 0.6125 ;
      RECT 94.27 0.3375 94.34 0.6125 ;
      RECT 94.485 0.2825 94.555 0.4175 ;
      RECT 94.27 0.3375 94.5575 0.4075 ;
      RECT 92.1775 1.455 93.305 1.525 ;
      RECT 93.235 0.725 93.305 1.525 ;
      RECT 92.1775 1.3125 92.2475 1.525 ;
      RECT 92.1475 1.3125 92.2825 1.3825 ;
      RECT 93.215 0.725 93.305 0.86 ;
      RECT 92.83 1.2375 92.9 1.3725 ;
      RECT 92.5175 1.2675 92.9 1.3375 ;
      RECT 92.44 0.8675 92.51 1.0025 ;
      RECT 92.29 0.8675 92.36 1.0025 ;
      RECT 91.855 0.8675 91.925 1.0025 ;
      RECT 91.515 0.8675 91.585 1.0025 ;
      RECT 91.515 0.9025 92.51 0.9725 ;
      RECT 91.675 0.6625 91.745 0.7975 ;
      RECT 91.135 0.6625 91.205 0.7975 ;
      RECT 91.135 0.695 91.745 0.765 ;
      RECT 90.895 0.87 90.965 1.005 ;
      RECT 90.755 0.87 90.825 1.005 ;
      RECT 91.335 0.8675 91.405 1.0025 ;
      RECT 90.755 0.9025 91.4075 0.9725 ;
      RECT 90.36 1.225 90.43 1.385 ;
      RECT 90.5925 1.225 90.7275 1.34 ;
      RECT 90.3625 0.5425 90.4325 1.32 ;
      RECT 90.36 1.225 90.7275 1.295 ;
      RECT 90.3625 0.5425 90.875 0.6125 ;
      RECT 90.805 0.3375 90.875 0.6125 ;
      RECT 91.02 0.2825 91.09 0.4175 ;
      RECT 90.805 0.3375 91.0925 0.4075 ;
      RECT 88.7125 1.455 89.84 1.525 ;
      RECT 89.77 0.725 89.84 1.525 ;
      RECT 88.7125 1.3125 88.7825 1.525 ;
      RECT 88.6825 1.3125 88.8175 1.3825 ;
      RECT 89.75 0.725 89.84 0.86 ;
      RECT 89.365 1.2375 89.435 1.3725 ;
      RECT 89.0525 1.2675 89.435 1.3375 ;
      RECT 88.975 0.8675 89.045 1.0025 ;
      RECT 88.825 0.8675 88.895 1.0025 ;
      RECT 88.39 0.8675 88.46 1.0025 ;
      RECT 88.05 0.8675 88.12 1.0025 ;
      RECT 88.05 0.9025 89.045 0.9725 ;
      RECT 88.21 0.6625 88.28 0.7975 ;
      RECT 87.67 0.6625 87.74 0.7975 ;
      RECT 87.67 0.695 88.28 0.765 ;
      RECT 87.43 0.87 87.5 1.005 ;
      RECT 87.29 0.87 87.36 1.005 ;
      RECT 87.87 0.8675 87.94 1.0025 ;
      RECT 87.29 0.9025 87.9425 0.9725 ;
      RECT 86.895 1.225 86.965 1.385 ;
      RECT 87.1275 1.225 87.2625 1.34 ;
      RECT 86.8975 0.5425 86.9675 1.32 ;
      RECT 86.895 1.225 87.2625 1.295 ;
      RECT 86.8975 0.5425 87.41 0.6125 ;
      RECT 87.34 0.3375 87.41 0.6125 ;
      RECT 87.555 0.2825 87.625 0.4175 ;
      RECT 87.34 0.3375 87.6275 0.4075 ;
      RECT 85.2475 1.455 86.375 1.525 ;
      RECT 86.305 0.725 86.375 1.525 ;
      RECT 85.2475 1.3125 85.3175 1.525 ;
      RECT 85.2175 1.3125 85.3525 1.3825 ;
      RECT 86.285 0.725 86.375 0.86 ;
      RECT 85.9 1.2375 85.97 1.3725 ;
      RECT 85.5875 1.2675 85.97 1.3375 ;
      RECT 85.51 0.8675 85.58 1.0025 ;
      RECT 85.36 0.8675 85.43 1.0025 ;
      RECT 84.925 0.8675 84.995 1.0025 ;
      RECT 84.585 0.8675 84.655 1.0025 ;
      RECT 84.585 0.9025 85.58 0.9725 ;
      RECT 84.745 0.6625 84.815 0.7975 ;
      RECT 84.205 0.6625 84.275 0.7975 ;
      RECT 84.205 0.695 84.815 0.765 ;
      RECT 83.965 0.87 84.035 1.005 ;
      RECT 83.825 0.87 83.895 1.005 ;
      RECT 84.405 0.8675 84.475 1.0025 ;
      RECT 83.825 0.9025 84.4775 0.9725 ;
      RECT 83.43 1.225 83.5 1.385 ;
      RECT 83.6625 1.225 83.7975 1.34 ;
      RECT 83.4325 0.5425 83.5025 1.32 ;
      RECT 83.43 1.225 83.7975 1.295 ;
      RECT 83.4325 0.5425 83.945 0.6125 ;
      RECT 83.875 0.3375 83.945 0.6125 ;
      RECT 84.09 0.2825 84.16 0.4175 ;
      RECT 83.875 0.3375 84.1625 0.4075 ;
      RECT 81.7825 1.455 82.91 1.525 ;
      RECT 82.84 0.725 82.91 1.525 ;
      RECT 81.7825 1.3125 81.8525 1.525 ;
      RECT 81.7525 1.3125 81.8875 1.3825 ;
      RECT 82.82 0.725 82.91 0.86 ;
      RECT 82.435 1.2375 82.505 1.3725 ;
      RECT 82.1225 1.2675 82.505 1.3375 ;
      RECT 82.045 0.8675 82.115 1.0025 ;
      RECT 81.895 0.8675 81.965 1.0025 ;
      RECT 81.46 0.8675 81.53 1.0025 ;
      RECT 81.12 0.8675 81.19 1.0025 ;
      RECT 81.12 0.9025 82.115 0.9725 ;
      RECT 81.28 0.6625 81.35 0.7975 ;
      RECT 80.74 0.6625 80.81 0.7975 ;
      RECT 80.74 0.695 81.35 0.765 ;
      RECT 80.5 0.87 80.57 1.005 ;
      RECT 80.36 0.87 80.43 1.005 ;
      RECT 80.94 0.8675 81.01 1.0025 ;
      RECT 80.36 0.9025 81.0125 0.9725 ;
      RECT 79.965 1.225 80.035 1.385 ;
      RECT 80.1975 1.225 80.3325 1.34 ;
      RECT 79.9675 0.5425 80.0375 1.32 ;
      RECT 79.965 1.225 80.3325 1.295 ;
      RECT 79.9675 0.5425 80.48 0.6125 ;
      RECT 80.41 0.3375 80.48 0.6125 ;
      RECT 80.625 0.2825 80.695 0.4175 ;
      RECT 80.41 0.3375 80.6975 0.4075 ;
      RECT 78.3175 1.455 79.445 1.525 ;
      RECT 79.375 0.725 79.445 1.525 ;
      RECT 78.3175 1.3125 78.3875 1.525 ;
      RECT 78.2875 1.3125 78.4225 1.3825 ;
      RECT 79.355 0.725 79.445 0.86 ;
      RECT 78.97 1.2375 79.04 1.3725 ;
      RECT 78.6575 1.2675 79.04 1.3375 ;
      RECT 78.58 0.8675 78.65 1.0025 ;
      RECT 78.43 0.8675 78.5 1.0025 ;
      RECT 77.995 0.8675 78.065 1.0025 ;
      RECT 77.655 0.8675 77.725 1.0025 ;
      RECT 77.655 0.9025 78.65 0.9725 ;
      RECT 77.815 0.6625 77.885 0.7975 ;
      RECT 77.275 0.6625 77.345 0.7975 ;
      RECT 77.275 0.695 77.885 0.765 ;
      RECT 77.035 0.87 77.105 1.005 ;
      RECT 76.895 0.87 76.965 1.005 ;
      RECT 77.475 0.8675 77.545 1.0025 ;
      RECT 76.895 0.9025 77.5475 0.9725 ;
      RECT 76.5 1.225 76.57 1.385 ;
      RECT 76.7325 1.225 76.8675 1.34 ;
      RECT 76.5025 0.5425 76.5725 1.32 ;
      RECT 76.5 1.225 76.8675 1.295 ;
      RECT 76.5025 0.5425 77.015 0.6125 ;
      RECT 76.945 0.3375 77.015 0.6125 ;
      RECT 77.16 0.2825 77.23 0.4175 ;
      RECT 76.945 0.3375 77.2325 0.4075 ;
      RECT 74.8525 1.455 75.98 1.525 ;
      RECT 75.91 0.725 75.98 1.525 ;
      RECT 74.8525 1.3125 74.9225 1.525 ;
      RECT 74.8225 1.3125 74.9575 1.3825 ;
      RECT 75.89 0.725 75.98 0.86 ;
      RECT 75.505 1.2375 75.575 1.3725 ;
      RECT 75.1925 1.2675 75.575 1.3375 ;
      RECT 75.115 0.8675 75.185 1.0025 ;
      RECT 74.965 0.8675 75.035 1.0025 ;
      RECT 74.53 0.8675 74.6 1.0025 ;
      RECT 74.19 0.8675 74.26 1.0025 ;
      RECT 74.19 0.9025 75.185 0.9725 ;
      RECT 74.35 0.6625 74.42 0.7975 ;
      RECT 73.81 0.6625 73.88 0.7975 ;
      RECT 73.81 0.695 74.42 0.765 ;
      RECT 73.57 0.87 73.64 1.005 ;
      RECT 73.43 0.87 73.5 1.005 ;
      RECT 74.01 0.8675 74.08 1.0025 ;
      RECT 73.43 0.9025 74.0825 0.9725 ;
      RECT 73.035 1.225 73.105 1.385 ;
      RECT 73.2675 1.225 73.4025 1.34 ;
      RECT 73.0375 0.5425 73.1075 1.32 ;
      RECT 73.035 1.225 73.4025 1.295 ;
      RECT 73.0375 0.5425 73.55 0.6125 ;
      RECT 73.48 0.3375 73.55 0.6125 ;
      RECT 73.695 0.2825 73.765 0.4175 ;
      RECT 73.48 0.3375 73.7675 0.4075 ;
      RECT 71.3875 1.455 72.515 1.525 ;
      RECT 72.445 0.725 72.515 1.525 ;
      RECT 71.3875 1.3125 71.4575 1.525 ;
      RECT 71.3575 1.3125 71.4925 1.3825 ;
      RECT 72.425 0.725 72.515 0.86 ;
      RECT 72.04 1.2375 72.11 1.3725 ;
      RECT 71.7275 1.2675 72.11 1.3375 ;
      RECT 71.65 0.8675 71.72 1.0025 ;
      RECT 71.5 0.8675 71.57 1.0025 ;
      RECT 71.065 0.8675 71.135 1.0025 ;
      RECT 70.725 0.8675 70.795 1.0025 ;
      RECT 70.725 0.9025 71.72 0.9725 ;
      RECT 70.885 0.6625 70.955 0.7975 ;
      RECT 70.345 0.6625 70.415 0.7975 ;
      RECT 70.345 0.695 70.955 0.765 ;
      RECT 70.105 0.87 70.175 1.005 ;
      RECT 69.965 0.87 70.035 1.005 ;
      RECT 70.545 0.8675 70.615 1.0025 ;
      RECT 69.965 0.9025 70.6175 0.9725 ;
      RECT 69.57 1.225 69.64 1.385 ;
      RECT 69.8025 1.225 69.9375 1.34 ;
      RECT 69.5725 0.5425 69.6425 1.32 ;
      RECT 69.57 1.225 69.9375 1.295 ;
      RECT 69.5725 0.5425 70.085 0.6125 ;
      RECT 70.015 0.3375 70.085 0.6125 ;
      RECT 70.23 0.2825 70.3 0.4175 ;
      RECT 70.015 0.3375 70.3025 0.4075 ;
      RECT 67.9225 1.455 69.05 1.525 ;
      RECT 68.98 0.725 69.05 1.525 ;
      RECT 67.9225 1.3125 67.9925 1.525 ;
      RECT 67.8925 1.3125 68.0275 1.3825 ;
      RECT 68.96 0.725 69.05 0.86 ;
      RECT 68.575 1.2375 68.645 1.3725 ;
      RECT 68.2625 1.2675 68.645 1.3375 ;
      RECT 68.185 0.8675 68.255 1.0025 ;
      RECT 68.035 0.8675 68.105 1.0025 ;
      RECT 67.6 0.8675 67.67 1.0025 ;
      RECT 67.26 0.8675 67.33 1.0025 ;
      RECT 67.26 0.9025 68.255 0.9725 ;
      RECT 67.42 0.6625 67.49 0.7975 ;
      RECT 66.88 0.6625 66.95 0.7975 ;
      RECT 66.88 0.695 67.49 0.765 ;
      RECT 66.64 0.87 66.71 1.005 ;
      RECT 66.5 0.87 66.57 1.005 ;
      RECT 67.08 0.8675 67.15 1.0025 ;
      RECT 66.5 0.9025 67.1525 0.9725 ;
      RECT 66.105 1.225 66.175 1.385 ;
      RECT 66.3375 1.225 66.4725 1.34 ;
      RECT 66.1075 0.5425 66.1775 1.32 ;
      RECT 66.105 1.225 66.4725 1.295 ;
      RECT 66.1075 0.5425 66.62 0.6125 ;
      RECT 66.55 0.3375 66.62 0.6125 ;
      RECT 66.765 0.2825 66.835 0.4175 ;
      RECT 66.55 0.3375 66.8375 0.4075 ;
      RECT 64.4575 1.455 65.585 1.525 ;
      RECT 65.515 0.725 65.585 1.525 ;
      RECT 64.4575 1.3125 64.5275 1.525 ;
      RECT 64.4275 1.3125 64.5625 1.3825 ;
      RECT 65.495 0.725 65.585 0.86 ;
      RECT 65.11 1.2375 65.18 1.3725 ;
      RECT 64.7975 1.2675 65.18 1.3375 ;
      RECT 64.72 0.8675 64.79 1.0025 ;
      RECT 64.57 0.8675 64.64 1.0025 ;
      RECT 64.135 0.8675 64.205 1.0025 ;
      RECT 63.795 0.8675 63.865 1.0025 ;
      RECT 63.795 0.9025 64.79 0.9725 ;
      RECT 63.955 0.6625 64.025 0.7975 ;
      RECT 63.415 0.6625 63.485 0.7975 ;
      RECT 63.415 0.695 64.025 0.765 ;
      RECT 63.175 0.87 63.245 1.005 ;
      RECT 63.035 0.87 63.105 1.005 ;
      RECT 63.615 0.8675 63.685 1.0025 ;
      RECT 63.035 0.9025 63.6875 0.9725 ;
      RECT 62.64 1.225 62.71 1.385 ;
      RECT 62.8725 1.225 63.0075 1.34 ;
      RECT 62.6425 0.5425 62.7125 1.32 ;
      RECT 62.64 1.225 63.0075 1.295 ;
      RECT 62.6425 0.5425 63.155 0.6125 ;
      RECT 63.085 0.3375 63.155 0.6125 ;
      RECT 63.3 0.2825 63.37 0.4175 ;
      RECT 63.085 0.3375 63.3725 0.4075 ;
      RECT 60.9925 1.455 62.12 1.525 ;
      RECT 62.05 0.725 62.12 1.525 ;
      RECT 60.9925 1.3125 61.0625 1.525 ;
      RECT 60.9625 1.3125 61.0975 1.3825 ;
      RECT 62.03 0.725 62.12 0.86 ;
      RECT 61.645 1.2375 61.715 1.3725 ;
      RECT 61.3325 1.2675 61.715 1.3375 ;
      RECT 61.255 0.8675 61.325 1.0025 ;
      RECT 61.105 0.8675 61.175 1.0025 ;
      RECT 60.67 0.8675 60.74 1.0025 ;
      RECT 60.33 0.8675 60.4 1.0025 ;
      RECT 60.33 0.9025 61.325 0.9725 ;
      RECT 60.49 0.6625 60.56 0.7975 ;
      RECT 59.95 0.6625 60.02 0.7975 ;
      RECT 59.95 0.695 60.56 0.765 ;
      RECT 59.71 0.87 59.78 1.005 ;
      RECT 59.57 0.87 59.64 1.005 ;
      RECT 60.15 0.8675 60.22 1.0025 ;
      RECT 59.57 0.9025 60.2225 0.9725 ;
      RECT 59.175 1.225 59.245 1.385 ;
      RECT 59.4075 1.225 59.5425 1.34 ;
      RECT 59.1775 0.5425 59.2475 1.32 ;
      RECT 59.175 1.225 59.5425 1.295 ;
      RECT 59.1775 0.5425 59.69 0.6125 ;
      RECT 59.62 0.3375 59.69 0.6125 ;
      RECT 59.835 0.2825 59.905 0.4175 ;
      RECT 59.62 0.3375 59.9075 0.4075 ;
      RECT 57.5275 1.455 58.655 1.525 ;
      RECT 58.585 0.725 58.655 1.525 ;
      RECT 57.5275 1.3125 57.5975 1.525 ;
      RECT 57.4975 1.3125 57.6325 1.3825 ;
      RECT 58.565 0.725 58.655 0.86 ;
      RECT 58.18 1.2375 58.25 1.3725 ;
      RECT 57.8675 1.2675 58.25 1.3375 ;
      RECT 57.79 0.8675 57.86 1.0025 ;
      RECT 57.64 0.8675 57.71 1.0025 ;
      RECT 57.205 0.8675 57.275 1.0025 ;
      RECT 56.865 0.8675 56.935 1.0025 ;
      RECT 56.865 0.9025 57.86 0.9725 ;
      RECT 57.025 0.6625 57.095 0.7975 ;
      RECT 56.485 0.6625 56.555 0.7975 ;
      RECT 56.485 0.695 57.095 0.765 ;
      RECT 56.245 0.87 56.315 1.005 ;
      RECT 56.105 0.87 56.175 1.005 ;
      RECT 56.685 0.8675 56.755 1.0025 ;
      RECT 56.105 0.9025 56.7575 0.9725 ;
      RECT 55.71 1.225 55.78 1.385 ;
      RECT 55.9425 1.225 56.0775 1.34 ;
      RECT 55.7125 0.5425 55.7825 1.32 ;
      RECT 55.71 1.225 56.0775 1.295 ;
      RECT 55.7125 0.5425 56.225 0.6125 ;
      RECT 56.155 0.3375 56.225 0.6125 ;
      RECT 56.37 0.2825 56.44 0.4175 ;
      RECT 56.155 0.3375 56.4425 0.4075 ;
      RECT 54.0625 1.455 55.19 1.525 ;
      RECT 55.12 0.725 55.19 1.525 ;
      RECT 54.0625 1.3125 54.1325 1.525 ;
      RECT 54.0325 1.3125 54.1675 1.3825 ;
      RECT 55.1 0.725 55.19 0.86 ;
      RECT 54.715 1.2375 54.785 1.3725 ;
      RECT 54.4025 1.2675 54.785 1.3375 ;
      RECT 54.325 0.8675 54.395 1.0025 ;
      RECT 54.175 0.8675 54.245 1.0025 ;
      RECT 53.74 0.8675 53.81 1.0025 ;
      RECT 53.4 0.8675 53.47 1.0025 ;
      RECT 53.4 0.9025 54.395 0.9725 ;
      RECT 53.56 0.6625 53.63 0.7975 ;
      RECT 53.02 0.6625 53.09 0.7975 ;
      RECT 53.02 0.695 53.63 0.765 ;
      RECT 52.78 0.87 52.85 1.005 ;
      RECT 52.64 0.87 52.71 1.005 ;
      RECT 53.22 0.8675 53.29 1.0025 ;
      RECT 52.64 0.9025 53.2925 0.9725 ;
      RECT 52.245 1.225 52.315 1.385 ;
      RECT 52.4775 1.225 52.6125 1.34 ;
      RECT 52.2475 0.5425 52.3175 1.32 ;
      RECT 52.245 1.225 52.6125 1.295 ;
      RECT 52.2475 0.5425 52.76 0.6125 ;
      RECT 52.69 0.3375 52.76 0.6125 ;
      RECT 52.905 0.2825 52.975 0.4175 ;
      RECT 52.69 0.3375 52.9775 0.4075 ;
      RECT 50.5975 1.455 51.725 1.525 ;
      RECT 51.655 0.725 51.725 1.525 ;
      RECT 50.5975 1.3125 50.6675 1.525 ;
      RECT 50.5675 1.3125 50.7025 1.3825 ;
      RECT 51.635 0.725 51.725 0.86 ;
      RECT 51.25 1.2375 51.32 1.3725 ;
      RECT 50.9375 1.2675 51.32 1.3375 ;
      RECT 50.86 0.8675 50.93 1.0025 ;
      RECT 50.71 0.8675 50.78 1.0025 ;
      RECT 50.275 0.8675 50.345 1.0025 ;
      RECT 49.935 0.8675 50.005 1.0025 ;
      RECT 49.935 0.9025 50.93 0.9725 ;
      RECT 50.095 0.6625 50.165 0.7975 ;
      RECT 49.555 0.6625 49.625 0.7975 ;
      RECT 49.555 0.695 50.165 0.765 ;
      RECT 49.315 0.87 49.385 1.005 ;
      RECT 49.175 0.87 49.245 1.005 ;
      RECT 49.755 0.8675 49.825 1.0025 ;
      RECT 49.175 0.9025 49.8275 0.9725 ;
      RECT 48.78 1.225 48.85 1.385 ;
      RECT 49.0125 1.225 49.1475 1.34 ;
      RECT 48.7825 0.5425 48.8525 1.32 ;
      RECT 48.78 1.225 49.1475 1.295 ;
      RECT 48.7825 0.5425 49.295 0.6125 ;
      RECT 49.225 0.3375 49.295 0.6125 ;
      RECT 49.44 0.2825 49.51 0.4175 ;
      RECT 49.225 0.3375 49.5125 0.4075 ;
      RECT 47.1325 1.455 48.26 1.525 ;
      RECT 48.19 0.725 48.26 1.525 ;
      RECT 47.1325 1.3125 47.2025 1.525 ;
      RECT 47.1025 1.3125 47.2375 1.3825 ;
      RECT 48.17 0.725 48.26 0.86 ;
      RECT 47.785 1.2375 47.855 1.3725 ;
      RECT 47.4725 1.2675 47.855 1.3375 ;
      RECT 47.395 0.8675 47.465 1.0025 ;
      RECT 47.245 0.8675 47.315 1.0025 ;
      RECT 46.81 0.8675 46.88 1.0025 ;
      RECT 46.47 0.8675 46.54 1.0025 ;
      RECT 46.47 0.9025 47.465 0.9725 ;
      RECT 46.63 0.6625 46.7 0.7975 ;
      RECT 46.09 0.6625 46.16 0.7975 ;
      RECT 46.09 0.695 46.7 0.765 ;
      RECT 45.85 0.87 45.92 1.005 ;
      RECT 45.71 0.87 45.78 1.005 ;
      RECT 46.29 0.8675 46.36 1.0025 ;
      RECT 45.71 0.9025 46.3625 0.9725 ;
      RECT 45.315 1.225 45.385 1.385 ;
      RECT 45.5475 1.225 45.6825 1.34 ;
      RECT 45.3175 0.5425 45.3875 1.32 ;
      RECT 45.315 1.225 45.6825 1.295 ;
      RECT 45.3175 0.5425 45.83 0.6125 ;
      RECT 45.76 0.3375 45.83 0.6125 ;
      RECT 45.975 0.2825 46.045 0.4175 ;
      RECT 45.76 0.3375 46.0475 0.4075 ;
      RECT 43.6675 1.455 44.795 1.525 ;
      RECT 44.725 0.725 44.795 1.525 ;
      RECT 43.6675 1.3125 43.7375 1.525 ;
      RECT 43.6375 1.3125 43.7725 1.3825 ;
      RECT 44.705 0.725 44.795 0.86 ;
      RECT 44.32 1.2375 44.39 1.3725 ;
      RECT 44.0075 1.2675 44.39 1.3375 ;
      RECT 43.93 0.8675 44 1.0025 ;
      RECT 43.78 0.8675 43.85 1.0025 ;
      RECT 43.345 0.8675 43.415 1.0025 ;
      RECT 43.005 0.8675 43.075 1.0025 ;
      RECT 43.005 0.9025 44 0.9725 ;
      RECT 43.165 0.6625 43.235 0.7975 ;
      RECT 42.625 0.6625 42.695 0.7975 ;
      RECT 42.625 0.695 43.235 0.765 ;
      RECT 42.385 0.87 42.455 1.005 ;
      RECT 42.245 0.87 42.315 1.005 ;
      RECT 42.825 0.8675 42.895 1.0025 ;
      RECT 42.245 0.9025 42.8975 0.9725 ;
      RECT 41.85 1.225 41.92 1.385 ;
      RECT 42.0825 1.225 42.2175 1.34 ;
      RECT 41.8525 0.5425 41.9225 1.32 ;
      RECT 41.85 1.225 42.2175 1.295 ;
      RECT 41.8525 0.5425 42.365 0.6125 ;
      RECT 42.295 0.3375 42.365 0.6125 ;
      RECT 42.51 0.2825 42.58 0.4175 ;
      RECT 42.295 0.3375 42.5825 0.4075 ;
      RECT 40.2025 1.455 41.33 1.525 ;
      RECT 41.26 0.725 41.33 1.525 ;
      RECT 40.2025 1.3125 40.2725 1.525 ;
      RECT 40.1725 1.3125 40.3075 1.3825 ;
      RECT 41.24 0.725 41.33 0.86 ;
      RECT 40.855 1.2375 40.925 1.3725 ;
      RECT 40.5425 1.2675 40.925 1.3375 ;
      RECT 40.465 0.8675 40.535 1.0025 ;
      RECT 40.315 0.8675 40.385 1.0025 ;
      RECT 39.88 0.8675 39.95 1.0025 ;
      RECT 39.54 0.8675 39.61 1.0025 ;
      RECT 39.54 0.9025 40.535 0.9725 ;
      RECT 39.7 0.6625 39.77 0.7975 ;
      RECT 39.16 0.6625 39.23 0.7975 ;
      RECT 39.16 0.695 39.77 0.765 ;
      RECT 38.92 0.87 38.99 1.005 ;
      RECT 38.78 0.87 38.85 1.005 ;
      RECT 39.36 0.8675 39.43 1.0025 ;
      RECT 38.78 0.9025 39.4325 0.9725 ;
      RECT 38.385 1.225 38.455 1.385 ;
      RECT 38.6175 1.225 38.7525 1.34 ;
      RECT 38.3875 0.5425 38.4575 1.32 ;
      RECT 38.385 1.225 38.7525 1.295 ;
      RECT 38.3875 0.5425 38.9 0.6125 ;
      RECT 38.83 0.3375 38.9 0.6125 ;
      RECT 39.045 0.2825 39.115 0.4175 ;
      RECT 38.83 0.3375 39.1175 0.4075 ;
      RECT 36.7375 1.455 37.865 1.525 ;
      RECT 37.795 0.725 37.865 1.525 ;
      RECT 36.7375 1.3125 36.8075 1.525 ;
      RECT 36.7075 1.3125 36.8425 1.3825 ;
      RECT 37.775 0.725 37.865 0.86 ;
      RECT 37.39 1.2375 37.46 1.3725 ;
      RECT 37.0775 1.2675 37.46 1.3375 ;
      RECT 37 0.8675 37.07 1.0025 ;
      RECT 36.85 0.8675 36.92 1.0025 ;
      RECT 36.415 0.8675 36.485 1.0025 ;
      RECT 36.075 0.8675 36.145 1.0025 ;
      RECT 36.075 0.9025 37.07 0.9725 ;
      RECT 36.235 0.6625 36.305 0.7975 ;
      RECT 35.695 0.6625 35.765 0.7975 ;
      RECT 35.695 0.695 36.305 0.765 ;
      RECT 35.455 0.87 35.525 1.005 ;
      RECT 35.315 0.87 35.385 1.005 ;
      RECT 35.895 0.8675 35.965 1.0025 ;
      RECT 35.315 0.9025 35.9675 0.9725 ;
      RECT 34.92 1.225 34.99 1.385 ;
      RECT 35.1525 1.225 35.2875 1.34 ;
      RECT 34.9225 0.5425 34.9925 1.32 ;
      RECT 34.92 1.225 35.2875 1.295 ;
      RECT 34.9225 0.5425 35.435 0.6125 ;
      RECT 35.365 0.3375 35.435 0.6125 ;
      RECT 35.58 0.2825 35.65 0.4175 ;
      RECT 35.365 0.3375 35.6525 0.4075 ;
      RECT 33.2725 1.455 34.4 1.525 ;
      RECT 34.33 0.725 34.4 1.525 ;
      RECT 33.2725 1.3125 33.3425 1.525 ;
      RECT 33.2425 1.3125 33.3775 1.3825 ;
      RECT 34.31 0.725 34.4 0.86 ;
      RECT 33.925 1.2375 33.995 1.3725 ;
      RECT 33.6125 1.2675 33.995 1.3375 ;
      RECT 33.535 0.8675 33.605 1.0025 ;
      RECT 33.385 0.8675 33.455 1.0025 ;
      RECT 32.95 0.8675 33.02 1.0025 ;
      RECT 32.61 0.8675 32.68 1.0025 ;
      RECT 32.61 0.9025 33.605 0.9725 ;
      RECT 32.77 0.6625 32.84 0.7975 ;
      RECT 32.23 0.6625 32.3 0.7975 ;
      RECT 32.23 0.695 32.84 0.765 ;
      RECT 31.99 0.87 32.06 1.005 ;
      RECT 31.85 0.87 31.92 1.005 ;
      RECT 32.43 0.8675 32.5 1.0025 ;
      RECT 31.85 0.9025 32.5025 0.9725 ;
      RECT 31.455 1.225 31.525 1.385 ;
      RECT 31.6875 1.225 31.8225 1.34 ;
      RECT 31.4575 0.5425 31.5275 1.32 ;
      RECT 31.455 1.225 31.8225 1.295 ;
      RECT 31.4575 0.5425 31.97 0.6125 ;
      RECT 31.9 0.3375 31.97 0.6125 ;
      RECT 32.115 0.2825 32.185 0.4175 ;
      RECT 31.9 0.3375 32.1875 0.4075 ;
      RECT 29.8075 1.455 30.935 1.525 ;
      RECT 30.865 0.725 30.935 1.525 ;
      RECT 29.8075 1.3125 29.8775 1.525 ;
      RECT 29.7775 1.3125 29.9125 1.3825 ;
      RECT 30.845 0.725 30.935 0.86 ;
      RECT 30.46 1.2375 30.53 1.3725 ;
      RECT 30.1475 1.2675 30.53 1.3375 ;
      RECT 30.07 0.8675 30.14 1.0025 ;
      RECT 29.92 0.8675 29.99 1.0025 ;
      RECT 29.485 0.8675 29.555 1.0025 ;
      RECT 29.145 0.8675 29.215 1.0025 ;
      RECT 29.145 0.9025 30.14 0.9725 ;
      RECT 29.305 0.6625 29.375 0.7975 ;
      RECT 28.765 0.6625 28.835 0.7975 ;
      RECT 28.765 0.695 29.375 0.765 ;
      RECT 28.525 0.87 28.595 1.005 ;
      RECT 28.385 0.87 28.455 1.005 ;
      RECT 28.965 0.8675 29.035 1.0025 ;
      RECT 28.385 0.9025 29.0375 0.9725 ;
      RECT 27.99 1.225 28.06 1.385 ;
      RECT 28.2225 1.225 28.3575 1.34 ;
      RECT 27.9925 0.5425 28.0625 1.32 ;
      RECT 27.99 1.225 28.3575 1.295 ;
      RECT 27.9925 0.5425 28.505 0.6125 ;
      RECT 28.435 0.3375 28.505 0.6125 ;
      RECT 28.65 0.2825 28.72 0.4175 ;
      RECT 28.435 0.3375 28.7225 0.4075 ;
      RECT 26.3425 1.455 27.47 1.525 ;
      RECT 27.4 0.725 27.47 1.525 ;
      RECT 26.3425 1.3125 26.4125 1.525 ;
      RECT 26.3125 1.3125 26.4475 1.3825 ;
      RECT 27.38 0.725 27.47 0.86 ;
      RECT 26.995 1.2375 27.065 1.3725 ;
      RECT 26.6825 1.2675 27.065 1.3375 ;
      RECT 26.605 0.8675 26.675 1.0025 ;
      RECT 26.455 0.8675 26.525 1.0025 ;
      RECT 26.02 0.8675 26.09 1.0025 ;
      RECT 25.68 0.8675 25.75 1.0025 ;
      RECT 25.68 0.9025 26.675 0.9725 ;
      RECT 25.84 0.6625 25.91 0.7975 ;
      RECT 25.3 0.6625 25.37 0.7975 ;
      RECT 25.3 0.695 25.91 0.765 ;
      RECT 25.06 0.87 25.13 1.005 ;
      RECT 24.92 0.87 24.99 1.005 ;
      RECT 25.5 0.8675 25.57 1.0025 ;
      RECT 24.92 0.9025 25.5725 0.9725 ;
      RECT 24.525 1.225 24.595 1.385 ;
      RECT 24.7575 1.225 24.8925 1.34 ;
      RECT 24.5275 0.5425 24.5975 1.32 ;
      RECT 24.525 1.225 24.8925 1.295 ;
      RECT 24.5275 0.5425 25.04 0.6125 ;
      RECT 24.97 0.3375 25.04 0.6125 ;
      RECT 25.185 0.2825 25.255 0.4175 ;
      RECT 24.97 0.3375 25.2575 0.4075 ;
      RECT 22.8775 1.455 24.005 1.525 ;
      RECT 23.935 0.725 24.005 1.525 ;
      RECT 22.8775 1.3125 22.9475 1.525 ;
      RECT 22.8475 1.3125 22.9825 1.3825 ;
      RECT 23.915 0.725 24.005 0.86 ;
      RECT 23.53 1.2375 23.6 1.3725 ;
      RECT 23.2175 1.2675 23.6 1.3375 ;
      RECT 23.14 0.8675 23.21 1.0025 ;
      RECT 22.99 0.8675 23.06 1.0025 ;
      RECT 22.555 0.8675 22.625 1.0025 ;
      RECT 22.215 0.8675 22.285 1.0025 ;
      RECT 22.215 0.9025 23.21 0.9725 ;
      RECT 22.375 0.6625 22.445 0.7975 ;
      RECT 21.835 0.6625 21.905 0.7975 ;
      RECT 21.835 0.695 22.445 0.765 ;
      RECT 21.595 0.87 21.665 1.005 ;
      RECT 21.455 0.87 21.525 1.005 ;
      RECT 22.035 0.8675 22.105 1.0025 ;
      RECT 21.455 0.9025 22.1075 0.9725 ;
      RECT 21.06 1.225 21.13 1.385 ;
      RECT 21.2925 1.225 21.4275 1.34 ;
      RECT 21.0625 0.5425 21.1325 1.32 ;
      RECT 21.06 1.225 21.4275 1.295 ;
      RECT 21.0625 0.5425 21.575 0.6125 ;
      RECT 21.505 0.3375 21.575 0.6125 ;
      RECT 21.72 0.2825 21.79 0.4175 ;
      RECT 21.505 0.3375 21.7925 0.4075 ;
      RECT 19.4125 1.455 20.54 1.525 ;
      RECT 20.47 0.725 20.54 1.525 ;
      RECT 19.4125 1.3125 19.4825 1.525 ;
      RECT 19.3825 1.3125 19.5175 1.3825 ;
      RECT 20.45 0.725 20.54 0.86 ;
      RECT 20.065 1.2375 20.135 1.3725 ;
      RECT 19.7525 1.2675 20.135 1.3375 ;
      RECT 19.675 0.8675 19.745 1.0025 ;
      RECT 19.525 0.8675 19.595 1.0025 ;
      RECT 19.09 0.8675 19.16 1.0025 ;
      RECT 18.75 0.8675 18.82 1.0025 ;
      RECT 18.75 0.9025 19.745 0.9725 ;
      RECT 18.91 0.6625 18.98 0.7975 ;
      RECT 18.37 0.6625 18.44 0.7975 ;
      RECT 18.37 0.695 18.98 0.765 ;
      RECT 18.13 0.87 18.2 1.005 ;
      RECT 17.99 0.87 18.06 1.005 ;
      RECT 18.57 0.8675 18.64 1.0025 ;
      RECT 17.99 0.9025 18.6425 0.9725 ;
      RECT 17.595 1.225 17.665 1.385 ;
      RECT 17.8275 1.225 17.9625 1.34 ;
      RECT 17.5975 0.5425 17.6675 1.32 ;
      RECT 17.595 1.225 17.9625 1.295 ;
      RECT 17.5975 0.5425 18.11 0.6125 ;
      RECT 18.04 0.3375 18.11 0.6125 ;
      RECT 18.255 0.2825 18.325 0.4175 ;
      RECT 18.04 0.3375 18.3275 0.4075 ;
      RECT 15.9475 1.455 17.075 1.525 ;
      RECT 17.005 0.725 17.075 1.525 ;
      RECT 15.9475 1.3125 16.0175 1.525 ;
      RECT 15.9175 1.3125 16.0525 1.3825 ;
      RECT 16.985 0.725 17.075 0.86 ;
      RECT 16.6 1.2375 16.67 1.3725 ;
      RECT 16.2875 1.2675 16.67 1.3375 ;
      RECT 16.21 0.8675 16.28 1.0025 ;
      RECT 16.06 0.8675 16.13 1.0025 ;
      RECT 15.625 0.8675 15.695 1.0025 ;
      RECT 15.285 0.8675 15.355 1.0025 ;
      RECT 15.285 0.9025 16.28 0.9725 ;
      RECT 15.445 0.6625 15.515 0.7975 ;
      RECT 14.905 0.6625 14.975 0.7975 ;
      RECT 14.905 0.695 15.515 0.765 ;
      RECT 14.665 0.87 14.735 1.005 ;
      RECT 14.525 0.87 14.595 1.005 ;
      RECT 15.105 0.8675 15.175 1.0025 ;
      RECT 14.525 0.9025 15.1775 0.9725 ;
      RECT 14.13 1.225 14.2 1.385 ;
      RECT 14.3625 1.225 14.4975 1.34 ;
      RECT 14.1325 0.5425 14.2025 1.32 ;
      RECT 14.13 1.225 14.4975 1.295 ;
      RECT 14.1325 0.5425 14.645 0.6125 ;
      RECT 14.575 0.3375 14.645 0.6125 ;
      RECT 14.79 0.2825 14.86 0.4175 ;
      RECT 14.575 0.3375 14.8625 0.4075 ;
      RECT 12.4825 1.455 13.61 1.525 ;
      RECT 13.54 0.725 13.61 1.525 ;
      RECT 12.4825 1.3125 12.5525 1.525 ;
      RECT 12.4525 1.3125 12.5875 1.3825 ;
      RECT 13.52 0.725 13.61 0.86 ;
      RECT 13.135 1.2375 13.205 1.3725 ;
      RECT 12.8225 1.2675 13.205 1.3375 ;
      RECT 12.745 0.8675 12.815 1.0025 ;
      RECT 12.595 0.8675 12.665 1.0025 ;
      RECT 12.16 0.8675 12.23 1.0025 ;
      RECT 11.82 0.8675 11.89 1.0025 ;
      RECT 11.82 0.9025 12.815 0.9725 ;
      RECT 11.98 0.6625 12.05 0.7975 ;
      RECT 11.44 0.6625 11.51 0.7975 ;
      RECT 11.44 0.695 12.05 0.765 ;
      RECT 11.2 0.87 11.27 1.005 ;
      RECT 11.06 0.87 11.13 1.005 ;
      RECT 11.64 0.8675 11.71 1.0025 ;
      RECT 11.06 0.9025 11.7125 0.9725 ;
      RECT 10.665 1.225 10.735 1.385 ;
      RECT 10.8975 1.225 11.0325 1.34 ;
      RECT 10.6675 0.5425 10.7375 1.32 ;
      RECT 10.665 1.225 11.0325 1.295 ;
      RECT 10.6675 0.5425 11.18 0.6125 ;
      RECT 11.11 0.3375 11.18 0.6125 ;
      RECT 11.325 0.2825 11.395 0.4175 ;
      RECT 11.11 0.3375 11.3975 0.4075 ;
      RECT 9.0175 1.455 10.145 1.525 ;
      RECT 10.075 0.725 10.145 1.525 ;
      RECT 9.0175 1.3125 9.0875 1.525 ;
      RECT 8.9875 1.3125 9.1225 1.3825 ;
      RECT 10.055 0.725 10.145 0.86 ;
      RECT 9.67 1.2375 9.74 1.3725 ;
      RECT 9.3575 1.2675 9.74 1.3375 ;
      RECT 9.28 0.8675 9.35 1.0025 ;
      RECT 9.13 0.8675 9.2 1.0025 ;
      RECT 8.695 0.8675 8.765 1.0025 ;
      RECT 8.355 0.8675 8.425 1.0025 ;
      RECT 8.355 0.9025 9.35 0.9725 ;
      RECT 8.515 0.6625 8.585 0.7975 ;
      RECT 7.975 0.6625 8.045 0.7975 ;
      RECT 7.975 0.695 8.585 0.765 ;
      RECT 7.735 0.87 7.805 1.005 ;
      RECT 7.595 0.87 7.665 1.005 ;
      RECT 8.175 0.8675 8.245 1.0025 ;
      RECT 7.595 0.9025 8.2475 0.9725 ;
      RECT 7.2 1.225 7.27 1.385 ;
      RECT 7.4325 1.225 7.5675 1.34 ;
      RECT 7.2025 0.5425 7.2725 1.32 ;
      RECT 7.2 1.225 7.5675 1.295 ;
      RECT 7.2025 0.5425 7.715 0.6125 ;
      RECT 7.645 0.3375 7.715 0.6125 ;
      RECT 7.86 0.2825 7.93 0.4175 ;
      RECT 7.645 0.3375 7.9325 0.4075 ;
      RECT 5.5525 1.455 6.68 1.525 ;
      RECT 6.61 0.725 6.68 1.525 ;
      RECT 5.5525 1.3125 5.6225 1.525 ;
      RECT 5.5225 1.3125 5.6575 1.3825 ;
      RECT 6.59 0.725 6.68 0.86 ;
      RECT 6.205 1.2375 6.275 1.3725 ;
      RECT 5.8925 1.2675 6.275 1.3375 ;
      RECT 5.815 0.8675 5.885 1.0025 ;
      RECT 5.665 0.8675 5.735 1.0025 ;
      RECT 5.23 0.8675 5.3 1.0025 ;
      RECT 4.89 0.8675 4.96 1.0025 ;
      RECT 4.89 0.9025 5.885 0.9725 ;
      RECT 5.05 0.6625 5.12 0.7975 ;
      RECT 4.51 0.6625 4.58 0.7975 ;
      RECT 4.51 0.695 5.12 0.765 ;
      RECT 4.27 0.87 4.34 1.005 ;
      RECT 4.13 0.87 4.2 1.005 ;
      RECT 4.71 0.8675 4.78 1.0025 ;
      RECT 4.13 0.9025 4.7825 0.9725 ;
      RECT 3.735 1.225 3.805 1.385 ;
      RECT 3.9675 1.225 4.1025 1.34 ;
      RECT 3.7375 0.5425 3.8075 1.32 ;
      RECT 3.735 1.225 4.1025 1.295 ;
      RECT 3.7375 0.5425 4.25 0.6125 ;
      RECT 4.18 0.3375 4.25 0.6125 ;
      RECT 4.395 0.2825 4.465 0.4175 ;
      RECT 4.18 0.3375 4.4675 0.4075 ;
      RECT 2.0875 1.455 3.215 1.525 ;
      RECT 3.145 0.725 3.215 1.525 ;
      RECT 2.0875 1.3125 2.1575 1.525 ;
      RECT 2.0575 1.3125 2.1925 1.3825 ;
      RECT 3.125 0.725 3.215 0.86 ;
      RECT 2.74 1.2375 2.81 1.3725 ;
      RECT 2.4275 1.2675 2.81 1.3375 ;
      RECT 2.35 0.8675 2.42 1.0025 ;
      RECT 2.2 0.8675 2.27 1.0025 ;
      RECT 1.765 0.8675 1.835 1.0025 ;
      RECT 1.425 0.8675 1.495 1.0025 ;
      RECT 1.425 0.9025 2.42 0.9725 ;
      RECT 1.585 0.6625 1.655 0.7975 ;
      RECT 1.045 0.6625 1.115 0.7975 ;
      RECT 1.045 0.695 1.655 0.765 ;
      RECT 0.805 0.87 0.875 1.005 ;
      RECT 0.665 0.87 0.735 1.005 ;
      RECT 1.245 0.8675 1.315 1.0025 ;
      RECT 0.665 0.9025 1.3175 0.9725 ;
      RECT 0.27 1.225 0.34 1.385 ;
      RECT 0.5025 1.225 0.6375 1.34 ;
      RECT 0.2725 0.5425 0.3425 1.32 ;
      RECT 0.27 1.225 0.6375 1.295 ;
      RECT 0.2725 0.5425 0.785 0.6125 ;
      RECT 0.715 0.3375 0.785 0.6125 ;
      RECT 0.93 0.2825 1 0.4175 ;
      RECT 0.715 0.3375 1.0025 0.4075 ;
      RECT 114.1325 0.705 114.2025 0.845 ;
      RECT 112.8825 0.45 112.9525 0.59 ;
      RECT 111.535 0.46 111.605 0.6 ;
      RECT 111.355 0.4525 111.425 0.5925 ;
      RECT 111.15 0.7175 111.22 0.8575 ;
      RECT 110.97 0.6775 111.04 0.8175 ;
      RECT 110.005 0.68 110.075 0.82 ;
      RECT 109.375 0.465 109.445 0.605 ;
      RECT 106.54 0.68 106.61 0.82 ;
      RECT 105.91 0.465 105.98 0.605 ;
      RECT 103.075 0.68 103.145 0.82 ;
      RECT 102.445 0.465 102.515 0.605 ;
      RECT 99.61 0.68 99.68 0.82 ;
      RECT 98.98 0.465 99.05 0.605 ;
      RECT 96.145 0.68 96.215 0.82 ;
      RECT 95.515 0.465 95.585 0.605 ;
      RECT 92.68 0.68 92.75 0.82 ;
      RECT 92.05 0.465 92.12 0.605 ;
      RECT 89.215 0.68 89.285 0.82 ;
      RECT 88.585 0.465 88.655 0.605 ;
      RECT 85.75 0.68 85.82 0.82 ;
      RECT 85.12 0.465 85.19 0.605 ;
      RECT 82.285 0.68 82.355 0.82 ;
      RECT 81.655 0.465 81.725 0.605 ;
      RECT 78.82 0.68 78.89 0.82 ;
      RECT 78.19 0.465 78.26 0.605 ;
      RECT 75.355 0.68 75.425 0.82 ;
      RECT 74.725 0.465 74.795 0.605 ;
      RECT 71.89 0.68 71.96 0.82 ;
      RECT 71.26 0.465 71.33 0.605 ;
      RECT 68.425 0.68 68.495 0.82 ;
      RECT 67.795 0.465 67.865 0.605 ;
      RECT 64.96 0.68 65.03 0.82 ;
      RECT 64.33 0.465 64.4 0.605 ;
      RECT 61.495 0.68 61.565 0.82 ;
      RECT 60.865 0.465 60.935 0.605 ;
      RECT 58.03 0.68 58.1 0.82 ;
      RECT 57.4 0.465 57.47 0.605 ;
      RECT 54.565 0.68 54.635 0.82 ;
      RECT 53.935 0.465 54.005 0.605 ;
      RECT 51.1 0.68 51.17 0.82 ;
      RECT 50.47 0.465 50.54 0.605 ;
      RECT 47.635 0.68 47.705 0.82 ;
      RECT 47.005 0.465 47.075 0.605 ;
      RECT 44.17 0.68 44.24 0.82 ;
      RECT 43.54 0.465 43.61 0.605 ;
      RECT 40.705 0.68 40.775 0.82 ;
      RECT 40.075 0.465 40.145 0.605 ;
      RECT 37.24 0.68 37.31 0.82 ;
      RECT 36.61 0.465 36.68 0.605 ;
      RECT 33.775 0.68 33.845 0.82 ;
      RECT 33.145 0.465 33.215 0.605 ;
      RECT 30.31 0.68 30.38 0.82 ;
      RECT 29.68 0.465 29.75 0.605 ;
      RECT 26.845 0.68 26.915 0.82 ;
      RECT 26.215 0.465 26.285 0.605 ;
      RECT 23.38 0.68 23.45 0.82 ;
      RECT 22.75 0.465 22.82 0.605 ;
      RECT 19.915 0.68 19.985 0.82 ;
      RECT 19.285 0.465 19.355 0.605 ;
      RECT 16.45 0.68 16.52 0.82 ;
      RECT 15.82 0.465 15.89 0.605 ;
      RECT 12.985 0.68 13.055 0.82 ;
      RECT 12.355 0.465 12.425 0.605 ;
      RECT 9.52 0.68 9.59 0.82 ;
      RECT 8.89 0.465 8.96 0.605 ;
      RECT 6.055 0.68 6.125 0.82 ;
      RECT 5.425 0.465 5.495 0.605 ;
      RECT 2.59 0.68 2.66 0.82 ;
      RECT 1.96 0.465 2.03 0.605 ;
    LAYER metal3 ;
      RECT 111.15 0.7175 111.22 0.8575 ;
      RECT 114.1325 0.705 114.2025 0.845 ;
      RECT 111.15 0.755 114.2025 0.825 ;
      RECT 111.535 0.46 111.605 0.6 ;
      RECT 112.8825 0.45 112.9525 0.59 ;
      RECT 111.535 0.4975 112.955 0.5675 ;
      RECT 109.375 0.125 109.445 0.605 ;
      RECT 105.91 0.125 105.98 0.605 ;
      RECT 102.445 0.125 102.515 0.605 ;
      RECT 98.98 0.125 99.05 0.605 ;
      RECT 95.515 0.125 95.585 0.605 ;
      RECT 92.05 0.125 92.12 0.605 ;
      RECT 88.585 0.125 88.655 0.605 ;
      RECT 85.12 0.125 85.19 0.605 ;
      RECT 81.655 0.125 81.725 0.605 ;
      RECT 78.19 0.125 78.26 0.605 ;
      RECT 74.725 0.125 74.795 0.605 ;
      RECT 71.26 0.125 71.33 0.605 ;
      RECT 67.795 0.125 67.865 0.605 ;
      RECT 64.33 0.125 64.4 0.605 ;
      RECT 60.865 0.125 60.935 0.605 ;
      RECT 57.4 0.125 57.47 0.605 ;
      RECT 53.935 0.125 54.005 0.605 ;
      RECT 50.47 0.125 50.54 0.605 ;
      RECT 47.005 0.125 47.075 0.605 ;
      RECT 43.54 0.125 43.61 0.605 ;
      RECT 40.075 0.125 40.145 0.605 ;
      RECT 36.61 0.125 36.68 0.605 ;
      RECT 33.145 0.125 33.215 0.605 ;
      RECT 29.68 0.125 29.75 0.605 ;
      RECT 26.215 0.125 26.285 0.605 ;
      RECT 22.75 0.125 22.82 0.605 ;
      RECT 19.285 0.125 19.355 0.605 ;
      RECT 15.82 0.125 15.89 0.605 ;
      RECT 12.355 0.125 12.425 0.605 ;
      RECT 8.89 0.125 8.96 0.605 ;
      RECT 5.425 0.125 5.495 0.605 ;
      RECT 1.96 0.125 2.03 0.605 ;
      RECT 111.355 0.4525 111.4275 0.5925 ;
      RECT 111.3575 0.125 111.4275 0.5925 ;
      RECT 1.96 0.125 111.4275 0.195 ;
      RECT 110.005 0.675 110.075 0.82 ;
      RECT 106.54 0.675 106.61 0.82 ;
      RECT 103.075 0.675 103.145 0.82 ;
      RECT 99.61 0.675 99.68 0.82 ;
      RECT 96.145 0.675 96.215 0.82 ;
      RECT 92.68 0.675 92.75 0.82 ;
      RECT 89.215 0.675 89.285 0.82 ;
      RECT 85.75 0.675 85.82 0.82 ;
      RECT 82.285 0.675 82.355 0.82 ;
      RECT 78.82 0.675 78.89 0.82 ;
      RECT 75.355 0.675 75.425 0.82 ;
      RECT 71.89 0.675 71.96 0.82 ;
      RECT 68.425 0.675 68.495 0.82 ;
      RECT 64.96 0.675 65.03 0.82 ;
      RECT 61.495 0.675 61.565 0.82 ;
      RECT 58.03 0.675 58.1 0.82 ;
      RECT 54.565 0.675 54.635 0.82 ;
      RECT 51.1 0.675 51.17 0.82 ;
      RECT 47.635 0.675 47.705 0.82 ;
      RECT 44.17 0.675 44.24 0.82 ;
      RECT 40.705 0.675 40.775 0.82 ;
      RECT 37.24 0.675 37.31 0.82 ;
      RECT 33.775 0.675 33.845 0.82 ;
      RECT 30.31 0.675 30.38 0.82 ;
      RECT 26.845 0.675 26.915 0.82 ;
      RECT 23.38 0.675 23.45 0.82 ;
      RECT 19.915 0.675 19.985 0.82 ;
      RECT 16.45 0.675 16.52 0.82 ;
      RECT 12.985 0.675 13.055 0.82 ;
      RECT 9.52 0.675 9.59 0.82 ;
      RECT 6.055 0.675 6.125 0.82 ;
      RECT 2.59 0.675 2.66 0.82 ;
      RECT 110.97 0.675 111.04 0.8175 ;
      RECT 2.59 0.675 111.0425 0.745 ;
    LAYER via1 ;
      RECT 115.17 1.065 115.235 1.13 ;
      RECT 114.715 0.44 114.78 0.505 ;
      RECT 114.715 0.995 114.78 1.06 ;
      RECT 114.585 1.255 114.65 1.32 ;
      RECT 114.455 0.44 114.52 0.505 ;
      RECT 114.455 1.05 114.52 1.115 ;
      RECT 114.135 0.7425 114.2 0.8075 ;
      RECT 113.98 0.5075 114.045 0.5725 ;
      RECT 113.98 1.2425 114.045 1.3075 ;
      RECT 113.7375 0.505 113.8025 0.57 ;
      RECT 113.6025 0.3 113.6675 0.365 ;
      RECT 113.4175 0.3 113.4825 0.365 ;
      RECT 113.2825 0.505 113.3475 0.57 ;
      RECT 113.04 0.5075 113.105 0.5725 ;
      RECT 113.04 1.2425 113.105 1.3075 ;
      RECT 112.885 0.4875 112.95 0.5525 ;
      RECT 112.565 0.44 112.63 0.505 ;
      RECT 112.565 1.05 112.63 1.115 ;
      RECT 112.435 1.255 112.5 1.32 ;
      RECT 112.305 0.44 112.37 0.505 ;
      RECT 112.305 0.995 112.37 1.06 ;
      RECT 111.85 1.065 111.915 1.13 ;
      RECT 111.5375 0.4975 111.6025 0.5625 ;
      RECT 111.3575 0.49 111.4225 0.555 ;
      RECT 111.1525 0.755 111.2175 0.82 ;
      RECT 110.9725 0.715 111.0375 0.78 ;
      RECT 110.5425 0.76 110.6075 0.825 ;
      RECT 110.1575 1.2725 110.2225 1.3375 ;
      RECT 110.0075 0.7175 110.0725 0.7825 ;
      RECT 109.8775 1.27 109.9425 1.335 ;
      RECT 109.7675 0.9025 109.8325 0.9675 ;
      RECT 109.6175 0.9025 109.6825 0.9675 ;
      RECT 109.5075 1.315 109.5725 1.38 ;
      RECT 109.3775 0.5025 109.4425 0.5675 ;
      RECT 109.1825 0.9025 109.2475 0.9675 ;
      RECT 109.0025 0.6975 109.0675 0.7625 ;
      RECT 108.8425 0.9025 108.9075 0.9675 ;
      RECT 108.6625 0.9025 108.7275 0.9675 ;
      RECT 108.4625 0.6975 108.5275 0.7625 ;
      RECT 108.3475 0.3175 108.4125 0.3825 ;
      RECT 108.2225 0.905 108.2875 0.97 ;
      RECT 108.0825 0.905 108.1475 0.97 ;
      RECT 107.9525 1.2725 108.0175 1.3375 ;
      RECT 107.6875 1.285 107.7525 1.35 ;
      RECT 107.0775 0.76 107.1425 0.825 ;
      RECT 106.6925 1.2725 106.7575 1.3375 ;
      RECT 106.5425 0.7175 106.6075 0.7825 ;
      RECT 106.4125 1.27 106.4775 1.335 ;
      RECT 106.3025 0.9025 106.3675 0.9675 ;
      RECT 106.1525 0.9025 106.2175 0.9675 ;
      RECT 106.0425 1.315 106.1075 1.38 ;
      RECT 105.9125 0.5025 105.9775 0.5675 ;
      RECT 105.7175 0.9025 105.7825 0.9675 ;
      RECT 105.5375 0.6975 105.6025 0.7625 ;
      RECT 105.3775 0.9025 105.4425 0.9675 ;
      RECT 105.1975 0.9025 105.2625 0.9675 ;
      RECT 104.9975 0.6975 105.0625 0.7625 ;
      RECT 104.8825 0.3175 104.9475 0.3825 ;
      RECT 104.7575 0.905 104.8225 0.97 ;
      RECT 104.6175 0.905 104.6825 0.97 ;
      RECT 104.4875 1.2725 104.5525 1.3375 ;
      RECT 104.2225 1.285 104.2875 1.35 ;
      RECT 103.6125 0.76 103.6775 0.825 ;
      RECT 103.2275 1.2725 103.2925 1.3375 ;
      RECT 103.0775 0.7175 103.1425 0.7825 ;
      RECT 102.9475 1.27 103.0125 1.335 ;
      RECT 102.8375 0.9025 102.9025 0.9675 ;
      RECT 102.6875 0.9025 102.7525 0.9675 ;
      RECT 102.5775 1.315 102.6425 1.38 ;
      RECT 102.4475 0.5025 102.5125 0.5675 ;
      RECT 102.2525 0.9025 102.3175 0.9675 ;
      RECT 102.0725 0.6975 102.1375 0.7625 ;
      RECT 101.9125 0.9025 101.9775 0.9675 ;
      RECT 101.7325 0.9025 101.7975 0.9675 ;
      RECT 101.5325 0.6975 101.5975 0.7625 ;
      RECT 101.4175 0.3175 101.4825 0.3825 ;
      RECT 101.2925 0.905 101.3575 0.97 ;
      RECT 101.1525 0.905 101.2175 0.97 ;
      RECT 101.0225 1.2725 101.0875 1.3375 ;
      RECT 100.7575 1.285 100.8225 1.35 ;
      RECT 100.1475 0.76 100.2125 0.825 ;
      RECT 99.7625 1.2725 99.8275 1.3375 ;
      RECT 99.6125 0.7175 99.6775 0.7825 ;
      RECT 99.4825 1.27 99.5475 1.335 ;
      RECT 99.3725 0.9025 99.4375 0.9675 ;
      RECT 99.2225 0.9025 99.2875 0.9675 ;
      RECT 99.1125 1.315 99.1775 1.38 ;
      RECT 98.9825 0.5025 99.0475 0.5675 ;
      RECT 98.7875 0.9025 98.8525 0.9675 ;
      RECT 98.6075 0.6975 98.6725 0.7625 ;
      RECT 98.4475 0.9025 98.5125 0.9675 ;
      RECT 98.2675 0.9025 98.3325 0.9675 ;
      RECT 98.0675 0.6975 98.1325 0.7625 ;
      RECT 97.9525 0.3175 98.0175 0.3825 ;
      RECT 97.8275 0.905 97.8925 0.97 ;
      RECT 97.6875 0.905 97.7525 0.97 ;
      RECT 97.5575 1.2725 97.6225 1.3375 ;
      RECT 97.2925 1.285 97.3575 1.35 ;
      RECT 96.6825 0.76 96.7475 0.825 ;
      RECT 96.2975 1.2725 96.3625 1.3375 ;
      RECT 96.1475 0.7175 96.2125 0.7825 ;
      RECT 96.0175 1.27 96.0825 1.335 ;
      RECT 95.9075 0.9025 95.9725 0.9675 ;
      RECT 95.7575 0.9025 95.8225 0.9675 ;
      RECT 95.6475 1.315 95.7125 1.38 ;
      RECT 95.5175 0.5025 95.5825 0.5675 ;
      RECT 95.3225 0.9025 95.3875 0.9675 ;
      RECT 95.1425 0.6975 95.2075 0.7625 ;
      RECT 94.9825 0.9025 95.0475 0.9675 ;
      RECT 94.8025 0.9025 94.8675 0.9675 ;
      RECT 94.6025 0.6975 94.6675 0.7625 ;
      RECT 94.4875 0.3175 94.5525 0.3825 ;
      RECT 94.3625 0.905 94.4275 0.97 ;
      RECT 94.2225 0.905 94.2875 0.97 ;
      RECT 94.0925 1.2725 94.1575 1.3375 ;
      RECT 93.8275 1.285 93.8925 1.35 ;
      RECT 93.2175 0.76 93.2825 0.825 ;
      RECT 92.8325 1.2725 92.8975 1.3375 ;
      RECT 92.6825 0.7175 92.7475 0.7825 ;
      RECT 92.5525 1.27 92.6175 1.335 ;
      RECT 92.4425 0.9025 92.5075 0.9675 ;
      RECT 92.2925 0.9025 92.3575 0.9675 ;
      RECT 92.1825 1.315 92.2475 1.38 ;
      RECT 92.0525 0.5025 92.1175 0.5675 ;
      RECT 91.8575 0.9025 91.9225 0.9675 ;
      RECT 91.6775 0.6975 91.7425 0.7625 ;
      RECT 91.5175 0.9025 91.5825 0.9675 ;
      RECT 91.3375 0.9025 91.4025 0.9675 ;
      RECT 91.1375 0.6975 91.2025 0.7625 ;
      RECT 91.0225 0.3175 91.0875 0.3825 ;
      RECT 90.8975 0.905 90.9625 0.97 ;
      RECT 90.7575 0.905 90.8225 0.97 ;
      RECT 90.6275 1.2725 90.6925 1.3375 ;
      RECT 90.3625 1.285 90.4275 1.35 ;
      RECT 89.7525 0.76 89.8175 0.825 ;
      RECT 89.3675 1.2725 89.4325 1.3375 ;
      RECT 89.2175 0.7175 89.2825 0.7825 ;
      RECT 89.0875 1.27 89.1525 1.335 ;
      RECT 88.9775 0.9025 89.0425 0.9675 ;
      RECT 88.8275 0.9025 88.8925 0.9675 ;
      RECT 88.7175 1.315 88.7825 1.38 ;
      RECT 88.5875 0.5025 88.6525 0.5675 ;
      RECT 88.3925 0.9025 88.4575 0.9675 ;
      RECT 88.2125 0.6975 88.2775 0.7625 ;
      RECT 88.0525 0.9025 88.1175 0.9675 ;
      RECT 87.8725 0.9025 87.9375 0.9675 ;
      RECT 87.6725 0.6975 87.7375 0.7625 ;
      RECT 87.5575 0.3175 87.6225 0.3825 ;
      RECT 87.4325 0.905 87.4975 0.97 ;
      RECT 87.2925 0.905 87.3575 0.97 ;
      RECT 87.1625 1.2725 87.2275 1.3375 ;
      RECT 86.8975 1.285 86.9625 1.35 ;
      RECT 86.2875 0.76 86.3525 0.825 ;
      RECT 85.9025 1.2725 85.9675 1.3375 ;
      RECT 85.7525 0.7175 85.8175 0.7825 ;
      RECT 85.6225 1.27 85.6875 1.335 ;
      RECT 85.5125 0.9025 85.5775 0.9675 ;
      RECT 85.3625 0.9025 85.4275 0.9675 ;
      RECT 85.2525 1.315 85.3175 1.38 ;
      RECT 85.1225 0.5025 85.1875 0.5675 ;
      RECT 84.9275 0.9025 84.9925 0.9675 ;
      RECT 84.7475 0.6975 84.8125 0.7625 ;
      RECT 84.5875 0.9025 84.6525 0.9675 ;
      RECT 84.4075 0.9025 84.4725 0.9675 ;
      RECT 84.2075 0.6975 84.2725 0.7625 ;
      RECT 84.0925 0.3175 84.1575 0.3825 ;
      RECT 83.9675 0.905 84.0325 0.97 ;
      RECT 83.8275 0.905 83.8925 0.97 ;
      RECT 83.6975 1.2725 83.7625 1.3375 ;
      RECT 83.4325 1.285 83.4975 1.35 ;
      RECT 82.8225 0.76 82.8875 0.825 ;
      RECT 82.4375 1.2725 82.5025 1.3375 ;
      RECT 82.2875 0.7175 82.3525 0.7825 ;
      RECT 82.1575 1.27 82.2225 1.335 ;
      RECT 82.0475 0.9025 82.1125 0.9675 ;
      RECT 81.8975 0.9025 81.9625 0.9675 ;
      RECT 81.7875 1.315 81.8525 1.38 ;
      RECT 81.6575 0.5025 81.7225 0.5675 ;
      RECT 81.4625 0.9025 81.5275 0.9675 ;
      RECT 81.2825 0.6975 81.3475 0.7625 ;
      RECT 81.1225 0.9025 81.1875 0.9675 ;
      RECT 80.9425 0.9025 81.0075 0.9675 ;
      RECT 80.7425 0.6975 80.8075 0.7625 ;
      RECT 80.6275 0.3175 80.6925 0.3825 ;
      RECT 80.5025 0.905 80.5675 0.97 ;
      RECT 80.3625 0.905 80.4275 0.97 ;
      RECT 80.2325 1.2725 80.2975 1.3375 ;
      RECT 79.9675 1.285 80.0325 1.35 ;
      RECT 79.3575 0.76 79.4225 0.825 ;
      RECT 78.9725 1.2725 79.0375 1.3375 ;
      RECT 78.8225 0.7175 78.8875 0.7825 ;
      RECT 78.6925 1.27 78.7575 1.335 ;
      RECT 78.5825 0.9025 78.6475 0.9675 ;
      RECT 78.4325 0.9025 78.4975 0.9675 ;
      RECT 78.3225 1.315 78.3875 1.38 ;
      RECT 78.1925 0.5025 78.2575 0.5675 ;
      RECT 77.9975 0.9025 78.0625 0.9675 ;
      RECT 77.8175 0.6975 77.8825 0.7625 ;
      RECT 77.6575 0.9025 77.7225 0.9675 ;
      RECT 77.4775 0.9025 77.5425 0.9675 ;
      RECT 77.2775 0.6975 77.3425 0.7625 ;
      RECT 77.1625 0.3175 77.2275 0.3825 ;
      RECT 77.0375 0.905 77.1025 0.97 ;
      RECT 76.8975 0.905 76.9625 0.97 ;
      RECT 76.7675 1.2725 76.8325 1.3375 ;
      RECT 76.5025 1.285 76.5675 1.35 ;
      RECT 75.8925 0.76 75.9575 0.825 ;
      RECT 75.5075 1.2725 75.5725 1.3375 ;
      RECT 75.3575 0.7175 75.4225 0.7825 ;
      RECT 75.2275 1.27 75.2925 1.335 ;
      RECT 75.1175 0.9025 75.1825 0.9675 ;
      RECT 74.9675 0.9025 75.0325 0.9675 ;
      RECT 74.8575 1.315 74.9225 1.38 ;
      RECT 74.7275 0.5025 74.7925 0.5675 ;
      RECT 74.5325 0.9025 74.5975 0.9675 ;
      RECT 74.3525 0.6975 74.4175 0.7625 ;
      RECT 74.1925 0.9025 74.2575 0.9675 ;
      RECT 74.0125 0.9025 74.0775 0.9675 ;
      RECT 73.8125 0.6975 73.8775 0.7625 ;
      RECT 73.6975 0.3175 73.7625 0.3825 ;
      RECT 73.5725 0.905 73.6375 0.97 ;
      RECT 73.4325 0.905 73.4975 0.97 ;
      RECT 73.3025 1.2725 73.3675 1.3375 ;
      RECT 73.0375 1.285 73.1025 1.35 ;
      RECT 72.4275 0.76 72.4925 0.825 ;
      RECT 72.0425 1.2725 72.1075 1.3375 ;
      RECT 71.8925 0.7175 71.9575 0.7825 ;
      RECT 71.7625 1.27 71.8275 1.335 ;
      RECT 71.6525 0.9025 71.7175 0.9675 ;
      RECT 71.5025 0.9025 71.5675 0.9675 ;
      RECT 71.3925 1.315 71.4575 1.38 ;
      RECT 71.2625 0.5025 71.3275 0.5675 ;
      RECT 71.0675 0.9025 71.1325 0.9675 ;
      RECT 70.8875 0.6975 70.9525 0.7625 ;
      RECT 70.7275 0.9025 70.7925 0.9675 ;
      RECT 70.5475 0.9025 70.6125 0.9675 ;
      RECT 70.3475 0.6975 70.4125 0.7625 ;
      RECT 70.2325 0.3175 70.2975 0.3825 ;
      RECT 70.1075 0.905 70.1725 0.97 ;
      RECT 69.9675 0.905 70.0325 0.97 ;
      RECT 69.8375 1.2725 69.9025 1.3375 ;
      RECT 69.5725 1.285 69.6375 1.35 ;
      RECT 68.9625 0.76 69.0275 0.825 ;
      RECT 68.5775 1.2725 68.6425 1.3375 ;
      RECT 68.4275 0.7175 68.4925 0.7825 ;
      RECT 68.2975 1.27 68.3625 1.335 ;
      RECT 68.1875 0.9025 68.2525 0.9675 ;
      RECT 68.0375 0.9025 68.1025 0.9675 ;
      RECT 67.9275 1.315 67.9925 1.38 ;
      RECT 67.7975 0.5025 67.8625 0.5675 ;
      RECT 67.6025 0.9025 67.6675 0.9675 ;
      RECT 67.4225 0.6975 67.4875 0.7625 ;
      RECT 67.2625 0.9025 67.3275 0.9675 ;
      RECT 67.0825 0.9025 67.1475 0.9675 ;
      RECT 66.8825 0.6975 66.9475 0.7625 ;
      RECT 66.7675 0.3175 66.8325 0.3825 ;
      RECT 66.6425 0.905 66.7075 0.97 ;
      RECT 66.5025 0.905 66.5675 0.97 ;
      RECT 66.3725 1.2725 66.4375 1.3375 ;
      RECT 66.1075 1.285 66.1725 1.35 ;
      RECT 65.4975 0.76 65.5625 0.825 ;
      RECT 65.1125 1.2725 65.1775 1.3375 ;
      RECT 64.9625 0.7175 65.0275 0.7825 ;
      RECT 64.8325 1.27 64.8975 1.335 ;
      RECT 64.7225 0.9025 64.7875 0.9675 ;
      RECT 64.5725 0.9025 64.6375 0.9675 ;
      RECT 64.4625 1.315 64.5275 1.38 ;
      RECT 64.3325 0.5025 64.3975 0.5675 ;
      RECT 64.1375 0.9025 64.2025 0.9675 ;
      RECT 63.9575 0.6975 64.0225 0.7625 ;
      RECT 63.7975 0.9025 63.8625 0.9675 ;
      RECT 63.6175 0.9025 63.6825 0.9675 ;
      RECT 63.4175 0.6975 63.4825 0.7625 ;
      RECT 63.3025 0.3175 63.3675 0.3825 ;
      RECT 63.1775 0.905 63.2425 0.97 ;
      RECT 63.0375 0.905 63.1025 0.97 ;
      RECT 62.9075 1.2725 62.9725 1.3375 ;
      RECT 62.6425 1.285 62.7075 1.35 ;
      RECT 62.0325 0.76 62.0975 0.825 ;
      RECT 61.6475 1.2725 61.7125 1.3375 ;
      RECT 61.4975 0.7175 61.5625 0.7825 ;
      RECT 61.3675 1.27 61.4325 1.335 ;
      RECT 61.2575 0.9025 61.3225 0.9675 ;
      RECT 61.1075 0.9025 61.1725 0.9675 ;
      RECT 60.9975 1.315 61.0625 1.38 ;
      RECT 60.8675 0.5025 60.9325 0.5675 ;
      RECT 60.6725 0.9025 60.7375 0.9675 ;
      RECT 60.4925 0.6975 60.5575 0.7625 ;
      RECT 60.3325 0.9025 60.3975 0.9675 ;
      RECT 60.1525 0.9025 60.2175 0.9675 ;
      RECT 59.9525 0.6975 60.0175 0.7625 ;
      RECT 59.8375 0.3175 59.9025 0.3825 ;
      RECT 59.7125 0.905 59.7775 0.97 ;
      RECT 59.5725 0.905 59.6375 0.97 ;
      RECT 59.4425 1.2725 59.5075 1.3375 ;
      RECT 59.1775 1.285 59.2425 1.35 ;
      RECT 58.5675 0.76 58.6325 0.825 ;
      RECT 58.1825 1.2725 58.2475 1.3375 ;
      RECT 58.0325 0.7175 58.0975 0.7825 ;
      RECT 57.9025 1.27 57.9675 1.335 ;
      RECT 57.7925 0.9025 57.8575 0.9675 ;
      RECT 57.6425 0.9025 57.7075 0.9675 ;
      RECT 57.5325 1.315 57.5975 1.38 ;
      RECT 57.4025 0.5025 57.4675 0.5675 ;
      RECT 57.2075 0.9025 57.2725 0.9675 ;
      RECT 57.0275 0.6975 57.0925 0.7625 ;
      RECT 56.8675 0.9025 56.9325 0.9675 ;
      RECT 56.6875 0.9025 56.7525 0.9675 ;
      RECT 56.4875 0.6975 56.5525 0.7625 ;
      RECT 56.3725 0.3175 56.4375 0.3825 ;
      RECT 56.2475 0.905 56.3125 0.97 ;
      RECT 56.1075 0.905 56.1725 0.97 ;
      RECT 55.9775 1.2725 56.0425 1.3375 ;
      RECT 55.7125 1.285 55.7775 1.35 ;
      RECT 55.1025 0.76 55.1675 0.825 ;
      RECT 54.7175 1.2725 54.7825 1.3375 ;
      RECT 54.5675 0.7175 54.6325 0.7825 ;
      RECT 54.4375 1.27 54.5025 1.335 ;
      RECT 54.3275 0.9025 54.3925 0.9675 ;
      RECT 54.1775 0.9025 54.2425 0.9675 ;
      RECT 54.0675 1.315 54.1325 1.38 ;
      RECT 53.9375 0.5025 54.0025 0.5675 ;
      RECT 53.7425 0.9025 53.8075 0.9675 ;
      RECT 53.5625 0.6975 53.6275 0.7625 ;
      RECT 53.4025 0.9025 53.4675 0.9675 ;
      RECT 53.2225 0.9025 53.2875 0.9675 ;
      RECT 53.0225 0.6975 53.0875 0.7625 ;
      RECT 52.9075 0.3175 52.9725 0.3825 ;
      RECT 52.7825 0.905 52.8475 0.97 ;
      RECT 52.6425 0.905 52.7075 0.97 ;
      RECT 52.5125 1.2725 52.5775 1.3375 ;
      RECT 52.2475 1.285 52.3125 1.35 ;
      RECT 51.6375 0.76 51.7025 0.825 ;
      RECT 51.2525 1.2725 51.3175 1.3375 ;
      RECT 51.1025 0.7175 51.1675 0.7825 ;
      RECT 50.9725 1.27 51.0375 1.335 ;
      RECT 50.8625 0.9025 50.9275 0.9675 ;
      RECT 50.7125 0.9025 50.7775 0.9675 ;
      RECT 50.6025 1.315 50.6675 1.38 ;
      RECT 50.4725 0.5025 50.5375 0.5675 ;
      RECT 50.2775 0.9025 50.3425 0.9675 ;
      RECT 50.0975 0.6975 50.1625 0.7625 ;
      RECT 49.9375 0.9025 50.0025 0.9675 ;
      RECT 49.7575 0.9025 49.8225 0.9675 ;
      RECT 49.5575 0.6975 49.6225 0.7625 ;
      RECT 49.4425 0.3175 49.5075 0.3825 ;
      RECT 49.3175 0.905 49.3825 0.97 ;
      RECT 49.1775 0.905 49.2425 0.97 ;
      RECT 49.0475 1.2725 49.1125 1.3375 ;
      RECT 48.7825 1.285 48.8475 1.35 ;
      RECT 48.1725 0.76 48.2375 0.825 ;
      RECT 47.7875 1.2725 47.8525 1.3375 ;
      RECT 47.6375 0.7175 47.7025 0.7825 ;
      RECT 47.5075 1.27 47.5725 1.335 ;
      RECT 47.3975 0.9025 47.4625 0.9675 ;
      RECT 47.2475 0.9025 47.3125 0.9675 ;
      RECT 47.1375 1.315 47.2025 1.38 ;
      RECT 47.0075 0.5025 47.0725 0.5675 ;
      RECT 46.8125 0.9025 46.8775 0.9675 ;
      RECT 46.6325 0.6975 46.6975 0.7625 ;
      RECT 46.4725 0.9025 46.5375 0.9675 ;
      RECT 46.2925 0.9025 46.3575 0.9675 ;
      RECT 46.0925 0.6975 46.1575 0.7625 ;
      RECT 45.9775 0.3175 46.0425 0.3825 ;
      RECT 45.8525 0.905 45.9175 0.97 ;
      RECT 45.7125 0.905 45.7775 0.97 ;
      RECT 45.5825 1.2725 45.6475 1.3375 ;
      RECT 45.3175 1.285 45.3825 1.35 ;
      RECT 44.7075 0.76 44.7725 0.825 ;
      RECT 44.3225 1.2725 44.3875 1.3375 ;
      RECT 44.1725 0.7175 44.2375 0.7825 ;
      RECT 44.0425 1.27 44.1075 1.335 ;
      RECT 43.9325 0.9025 43.9975 0.9675 ;
      RECT 43.7825 0.9025 43.8475 0.9675 ;
      RECT 43.6725 1.315 43.7375 1.38 ;
      RECT 43.5425 0.5025 43.6075 0.5675 ;
      RECT 43.3475 0.9025 43.4125 0.9675 ;
      RECT 43.1675 0.6975 43.2325 0.7625 ;
      RECT 43.0075 0.9025 43.0725 0.9675 ;
      RECT 42.8275 0.9025 42.8925 0.9675 ;
      RECT 42.6275 0.6975 42.6925 0.7625 ;
      RECT 42.5125 0.3175 42.5775 0.3825 ;
      RECT 42.3875 0.905 42.4525 0.97 ;
      RECT 42.2475 0.905 42.3125 0.97 ;
      RECT 42.1175 1.2725 42.1825 1.3375 ;
      RECT 41.8525 1.285 41.9175 1.35 ;
      RECT 41.2425 0.76 41.3075 0.825 ;
      RECT 40.8575 1.2725 40.9225 1.3375 ;
      RECT 40.7075 0.7175 40.7725 0.7825 ;
      RECT 40.5775 1.27 40.6425 1.335 ;
      RECT 40.4675 0.9025 40.5325 0.9675 ;
      RECT 40.3175 0.9025 40.3825 0.9675 ;
      RECT 40.2075 1.315 40.2725 1.38 ;
      RECT 40.0775 0.5025 40.1425 0.5675 ;
      RECT 39.8825 0.9025 39.9475 0.9675 ;
      RECT 39.7025 0.6975 39.7675 0.7625 ;
      RECT 39.5425 0.9025 39.6075 0.9675 ;
      RECT 39.3625 0.9025 39.4275 0.9675 ;
      RECT 39.1625 0.6975 39.2275 0.7625 ;
      RECT 39.0475 0.3175 39.1125 0.3825 ;
      RECT 38.9225 0.905 38.9875 0.97 ;
      RECT 38.7825 0.905 38.8475 0.97 ;
      RECT 38.6525 1.2725 38.7175 1.3375 ;
      RECT 38.3875 1.285 38.4525 1.35 ;
      RECT 37.7775 0.76 37.8425 0.825 ;
      RECT 37.3925 1.2725 37.4575 1.3375 ;
      RECT 37.2425 0.7175 37.3075 0.7825 ;
      RECT 37.1125 1.27 37.1775 1.335 ;
      RECT 37.0025 0.9025 37.0675 0.9675 ;
      RECT 36.8525 0.9025 36.9175 0.9675 ;
      RECT 36.7425 1.315 36.8075 1.38 ;
      RECT 36.6125 0.5025 36.6775 0.5675 ;
      RECT 36.4175 0.9025 36.4825 0.9675 ;
      RECT 36.2375 0.6975 36.3025 0.7625 ;
      RECT 36.0775 0.9025 36.1425 0.9675 ;
      RECT 35.8975 0.9025 35.9625 0.9675 ;
      RECT 35.6975 0.6975 35.7625 0.7625 ;
      RECT 35.5825 0.3175 35.6475 0.3825 ;
      RECT 35.4575 0.905 35.5225 0.97 ;
      RECT 35.3175 0.905 35.3825 0.97 ;
      RECT 35.1875 1.2725 35.2525 1.3375 ;
      RECT 34.9225 1.285 34.9875 1.35 ;
      RECT 34.3125 0.76 34.3775 0.825 ;
      RECT 33.9275 1.2725 33.9925 1.3375 ;
      RECT 33.7775 0.7175 33.8425 0.7825 ;
      RECT 33.6475 1.27 33.7125 1.335 ;
      RECT 33.5375 0.9025 33.6025 0.9675 ;
      RECT 33.3875 0.9025 33.4525 0.9675 ;
      RECT 33.2775 1.315 33.3425 1.38 ;
      RECT 33.1475 0.5025 33.2125 0.5675 ;
      RECT 32.9525 0.9025 33.0175 0.9675 ;
      RECT 32.7725 0.6975 32.8375 0.7625 ;
      RECT 32.6125 0.9025 32.6775 0.9675 ;
      RECT 32.4325 0.9025 32.4975 0.9675 ;
      RECT 32.2325 0.6975 32.2975 0.7625 ;
      RECT 32.1175 0.3175 32.1825 0.3825 ;
      RECT 31.9925 0.905 32.0575 0.97 ;
      RECT 31.8525 0.905 31.9175 0.97 ;
      RECT 31.7225 1.2725 31.7875 1.3375 ;
      RECT 31.4575 1.285 31.5225 1.35 ;
      RECT 30.8475 0.76 30.9125 0.825 ;
      RECT 30.4625 1.2725 30.5275 1.3375 ;
      RECT 30.3125 0.7175 30.3775 0.7825 ;
      RECT 30.1825 1.27 30.2475 1.335 ;
      RECT 30.0725 0.9025 30.1375 0.9675 ;
      RECT 29.9225 0.9025 29.9875 0.9675 ;
      RECT 29.8125 1.315 29.8775 1.38 ;
      RECT 29.6825 0.5025 29.7475 0.5675 ;
      RECT 29.4875 0.9025 29.5525 0.9675 ;
      RECT 29.3075 0.6975 29.3725 0.7625 ;
      RECT 29.1475 0.9025 29.2125 0.9675 ;
      RECT 28.9675 0.9025 29.0325 0.9675 ;
      RECT 28.7675 0.6975 28.8325 0.7625 ;
      RECT 28.6525 0.3175 28.7175 0.3825 ;
      RECT 28.5275 0.905 28.5925 0.97 ;
      RECT 28.3875 0.905 28.4525 0.97 ;
      RECT 28.2575 1.2725 28.3225 1.3375 ;
      RECT 27.9925 1.285 28.0575 1.35 ;
      RECT 27.3825 0.76 27.4475 0.825 ;
      RECT 26.9975 1.2725 27.0625 1.3375 ;
      RECT 26.8475 0.7175 26.9125 0.7825 ;
      RECT 26.7175 1.27 26.7825 1.335 ;
      RECT 26.6075 0.9025 26.6725 0.9675 ;
      RECT 26.4575 0.9025 26.5225 0.9675 ;
      RECT 26.3475 1.315 26.4125 1.38 ;
      RECT 26.2175 0.5025 26.2825 0.5675 ;
      RECT 26.0225 0.9025 26.0875 0.9675 ;
      RECT 25.8425 0.6975 25.9075 0.7625 ;
      RECT 25.6825 0.9025 25.7475 0.9675 ;
      RECT 25.5025 0.9025 25.5675 0.9675 ;
      RECT 25.3025 0.6975 25.3675 0.7625 ;
      RECT 25.1875 0.3175 25.2525 0.3825 ;
      RECT 25.0625 0.905 25.1275 0.97 ;
      RECT 24.9225 0.905 24.9875 0.97 ;
      RECT 24.7925 1.2725 24.8575 1.3375 ;
      RECT 24.5275 1.285 24.5925 1.35 ;
      RECT 23.9175 0.76 23.9825 0.825 ;
      RECT 23.5325 1.2725 23.5975 1.3375 ;
      RECT 23.3825 0.7175 23.4475 0.7825 ;
      RECT 23.2525 1.27 23.3175 1.335 ;
      RECT 23.1425 0.9025 23.2075 0.9675 ;
      RECT 22.9925 0.9025 23.0575 0.9675 ;
      RECT 22.8825 1.315 22.9475 1.38 ;
      RECT 22.7525 0.5025 22.8175 0.5675 ;
      RECT 22.5575 0.9025 22.6225 0.9675 ;
      RECT 22.3775 0.6975 22.4425 0.7625 ;
      RECT 22.2175 0.9025 22.2825 0.9675 ;
      RECT 22.0375 0.9025 22.1025 0.9675 ;
      RECT 21.8375 0.6975 21.9025 0.7625 ;
      RECT 21.7225 0.3175 21.7875 0.3825 ;
      RECT 21.5975 0.905 21.6625 0.97 ;
      RECT 21.4575 0.905 21.5225 0.97 ;
      RECT 21.3275 1.2725 21.3925 1.3375 ;
      RECT 21.0625 1.285 21.1275 1.35 ;
      RECT 20.4525 0.76 20.5175 0.825 ;
      RECT 20.0675 1.2725 20.1325 1.3375 ;
      RECT 19.9175 0.7175 19.9825 0.7825 ;
      RECT 19.7875 1.27 19.8525 1.335 ;
      RECT 19.6775 0.9025 19.7425 0.9675 ;
      RECT 19.5275 0.9025 19.5925 0.9675 ;
      RECT 19.4175 1.315 19.4825 1.38 ;
      RECT 19.2875 0.5025 19.3525 0.5675 ;
      RECT 19.0925 0.9025 19.1575 0.9675 ;
      RECT 18.9125 0.6975 18.9775 0.7625 ;
      RECT 18.7525 0.9025 18.8175 0.9675 ;
      RECT 18.5725 0.9025 18.6375 0.9675 ;
      RECT 18.3725 0.6975 18.4375 0.7625 ;
      RECT 18.2575 0.3175 18.3225 0.3825 ;
      RECT 18.1325 0.905 18.1975 0.97 ;
      RECT 17.9925 0.905 18.0575 0.97 ;
      RECT 17.8625 1.2725 17.9275 1.3375 ;
      RECT 17.5975 1.285 17.6625 1.35 ;
      RECT 16.9875 0.76 17.0525 0.825 ;
      RECT 16.6025 1.2725 16.6675 1.3375 ;
      RECT 16.4525 0.7175 16.5175 0.7825 ;
      RECT 16.3225 1.27 16.3875 1.335 ;
      RECT 16.2125 0.9025 16.2775 0.9675 ;
      RECT 16.0625 0.9025 16.1275 0.9675 ;
      RECT 15.9525 1.315 16.0175 1.38 ;
      RECT 15.8225 0.5025 15.8875 0.5675 ;
      RECT 15.6275 0.9025 15.6925 0.9675 ;
      RECT 15.4475 0.6975 15.5125 0.7625 ;
      RECT 15.2875 0.9025 15.3525 0.9675 ;
      RECT 15.1075 0.9025 15.1725 0.9675 ;
      RECT 14.9075 0.6975 14.9725 0.7625 ;
      RECT 14.7925 0.3175 14.8575 0.3825 ;
      RECT 14.6675 0.905 14.7325 0.97 ;
      RECT 14.5275 0.905 14.5925 0.97 ;
      RECT 14.3975 1.2725 14.4625 1.3375 ;
      RECT 14.1325 1.285 14.1975 1.35 ;
      RECT 13.5225 0.76 13.5875 0.825 ;
      RECT 13.1375 1.2725 13.2025 1.3375 ;
      RECT 12.9875 0.7175 13.0525 0.7825 ;
      RECT 12.8575 1.27 12.9225 1.335 ;
      RECT 12.7475 0.9025 12.8125 0.9675 ;
      RECT 12.5975 0.9025 12.6625 0.9675 ;
      RECT 12.4875 1.315 12.5525 1.38 ;
      RECT 12.3575 0.5025 12.4225 0.5675 ;
      RECT 12.1625 0.9025 12.2275 0.9675 ;
      RECT 11.9825 0.6975 12.0475 0.7625 ;
      RECT 11.8225 0.9025 11.8875 0.9675 ;
      RECT 11.6425 0.9025 11.7075 0.9675 ;
      RECT 11.4425 0.6975 11.5075 0.7625 ;
      RECT 11.3275 0.3175 11.3925 0.3825 ;
      RECT 11.2025 0.905 11.2675 0.97 ;
      RECT 11.0625 0.905 11.1275 0.97 ;
      RECT 10.9325 1.2725 10.9975 1.3375 ;
      RECT 10.6675 1.285 10.7325 1.35 ;
      RECT 10.0575 0.76 10.1225 0.825 ;
      RECT 9.6725 1.2725 9.7375 1.3375 ;
      RECT 9.5225 0.7175 9.5875 0.7825 ;
      RECT 9.3925 1.27 9.4575 1.335 ;
      RECT 9.2825 0.9025 9.3475 0.9675 ;
      RECT 9.1325 0.9025 9.1975 0.9675 ;
      RECT 9.0225 1.315 9.0875 1.38 ;
      RECT 8.8925 0.5025 8.9575 0.5675 ;
      RECT 8.6975 0.9025 8.7625 0.9675 ;
      RECT 8.5175 0.6975 8.5825 0.7625 ;
      RECT 8.3575 0.9025 8.4225 0.9675 ;
      RECT 8.1775 0.9025 8.2425 0.9675 ;
      RECT 7.9775 0.6975 8.0425 0.7625 ;
      RECT 7.8625 0.3175 7.9275 0.3825 ;
      RECT 7.7375 0.905 7.8025 0.97 ;
      RECT 7.5975 0.905 7.6625 0.97 ;
      RECT 7.4675 1.2725 7.5325 1.3375 ;
      RECT 7.2025 1.285 7.2675 1.35 ;
      RECT 6.5925 0.76 6.6575 0.825 ;
      RECT 6.2075 1.2725 6.2725 1.3375 ;
      RECT 6.0575 0.7175 6.1225 0.7825 ;
      RECT 5.9275 1.27 5.9925 1.335 ;
      RECT 5.8175 0.9025 5.8825 0.9675 ;
      RECT 5.6675 0.9025 5.7325 0.9675 ;
      RECT 5.5575 1.315 5.6225 1.38 ;
      RECT 5.4275 0.5025 5.4925 0.5675 ;
      RECT 5.2325 0.9025 5.2975 0.9675 ;
      RECT 5.0525 0.6975 5.1175 0.7625 ;
      RECT 4.8925 0.9025 4.9575 0.9675 ;
      RECT 4.7125 0.9025 4.7775 0.9675 ;
      RECT 4.5125 0.6975 4.5775 0.7625 ;
      RECT 4.3975 0.3175 4.4625 0.3825 ;
      RECT 4.2725 0.905 4.3375 0.97 ;
      RECT 4.1325 0.905 4.1975 0.97 ;
      RECT 4.0025 1.2725 4.0675 1.3375 ;
      RECT 3.7375 1.285 3.8025 1.35 ;
      RECT 3.1275 0.76 3.1925 0.825 ;
      RECT 2.7425 1.2725 2.8075 1.3375 ;
      RECT 2.5925 0.7175 2.6575 0.7825 ;
      RECT 2.4625 1.27 2.5275 1.335 ;
      RECT 2.3525 0.9025 2.4175 0.9675 ;
      RECT 2.2025 0.9025 2.2675 0.9675 ;
      RECT 2.0925 1.315 2.1575 1.38 ;
      RECT 1.9625 0.5025 2.0275 0.5675 ;
      RECT 1.7675 0.9025 1.8325 0.9675 ;
      RECT 1.5875 0.6975 1.6525 0.7625 ;
      RECT 1.4275 0.9025 1.4925 0.9675 ;
      RECT 1.2475 0.9025 1.3125 0.9675 ;
      RECT 1.0475 0.6975 1.1125 0.7625 ;
      RECT 0.9325 0.3175 0.9975 0.3825 ;
      RECT 0.8075 0.905 0.8725 0.97 ;
      RECT 0.6675 0.905 0.7325 0.97 ;
      RECT 0.5375 1.2725 0.6025 1.3375 ;
      RECT 0.2725 1.285 0.3375 1.35 ;
    LAYER via2 ;
      RECT 114.1325 0.74 114.2025 0.81 ;
      RECT 112.8825 0.485 112.9525 0.555 ;
      RECT 111.535 0.495 111.605 0.565 ;
      RECT 111.355 0.4875 111.425 0.5575 ;
      RECT 111.15 0.7525 111.22 0.8225 ;
      RECT 110.97 0.7125 111.04 0.7825 ;
      RECT 110.005 0.715 110.075 0.785 ;
      RECT 109.375 0.5 109.445 0.57 ;
      RECT 106.54 0.715 106.61 0.785 ;
      RECT 105.91 0.5 105.98 0.57 ;
      RECT 103.075 0.715 103.145 0.785 ;
      RECT 102.445 0.5 102.515 0.57 ;
      RECT 99.61 0.715 99.68 0.785 ;
      RECT 98.98 0.5 99.05 0.57 ;
      RECT 96.145 0.715 96.215 0.785 ;
      RECT 95.515 0.5 95.585 0.57 ;
      RECT 92.68 0.715 92.75 0.785 ;
      RECT 92.05 0.5 92.12 0.57 ;
      RECT 89.215 0.715 89.285 0.785 ;
      RECT 88.585 0.5 88.655 0.57 ;
      RECT 85.75 0.715 85.82 0.785 ;
      RECT 85.12 0.5 85.19 0.57 ;
      RECT 82.285 0.715 82.355 0.785 ;
      RECT 81.655 0.5 81.725 0.57 ;
      RECT 78.82 0.715 78.89 0.785 ;
      RECT 78.19 0.5 78.26 0.57 ;
      RECT 75.355 0.715 75.425 0.785 ;
      RECT 74.725 0.5 74.795 0.57 ;
      RECT 71.89 0.715 71.96 0.785 ;
      RECT 71.26 0.5 71.33 0.57 ;
      RECT 68.425 0.715 68.495 0.785 ;
      RECT 67.795 0.5 67.865 0.57 ;
      RECT 64.96 0.715 65.03 0.785 ;
      RECT 64.33 0.5 64.4 0.57 ;
      RECT 61.495 0.715 61.565 0.785 ;
      RECT 60.865 0.5 60.935 0.57 ;
      RECT 58.03 0.715 58.1 0.785 ;
      RECT 57.4 0.5 57.47 0.57 ;
      RECT 54.565 0.715 54.635 0.785 ;
      RECT 53.935 0.5 54.005 0.57 ;
      RECT 51.1 0.715 51.17 0.785 ;
      RECT 50.47 0.5 50.54 0.57 ;
      RECT 47.635 0.715 47.705 0.785 ;
      RECT 47.005 0.5 47.075 0.57 ;
      RECT 44.17 0.715 44.24 0.785 ;
      RECT 43.54 0.5 43.61 0.57 ;
      RECT 40.705 0.715 40.775 0.785 ;
      RECT 40.075 0.5 40.145 0.57 ;
      RECT 37.24 0.715 37.31 0.785 ;
      RECT 36.61 0.5 36.68 0.57 ;
      RECT 33.775 0.715 33.845 0.785 ;
      RECT 33.145 0.5 33.215 0.57 ;
      RECT 30.31 0.715 30.38 0.785 ;
      RECT 29.68 0.5 29.75 0.57 ;
      RECT 26.845 0.715 26.915 0.785 ;
      RECT 26.215 0.5 26.285 0.57 ;
      RECT 23.38 0.715 23.45 0.785 ;
      RECT 22.75 0.5 22.82 0.57 ;
      RECT 19.915 0.715 19.985 0.785 ;
      RECT 19.285 0.5 19.355 0.57 ;
      RECT 16.45 0.715 16.52 0.785 ;
      RECT 15.82 0.5 15.89 0.57 ;
      RECT 12.985 0.715 13.055 0.785 ;
      RECT 12.355 0.5 12.425 0.57 ;
      RECT 9.52 0.715 9.59 0.785 ;
      RECT 8.89 0.5 8.96 0.57 ;
      RECT 6.055 0.715 6.125 0.785 ;
      RECT 5.425 0.5 5.495 0.57 ;
      RECT 2.59 0.715 2.66 0.785 ;
      RECT 1.96 0.5 2.03 0.57 ;
  END
END regfile

END LIBRARY
